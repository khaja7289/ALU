magic
tech scmos
timestamp 1696145522
<< metal1 >>
rect 992 3303 994 3307
rect 998 3303 1001 3307
rect 1005 3303 1008 3307
rect 2024 3303 2026 3307
rect 2030 3303 2033 3307
rect 2037 3303 2040 3307
rect 3040 3303 3042 3307
rect 3046 3303 3049 3307
rect 3053 3303 3056 3307
rect 494 3288 502 3291
rect 2394 3288 2395 3292
rect 2542 3288 2558 3291
rect 3046 3288 3062 3291
rect 150 3278 169 3281
rect 438 3278 449 3281
rect 366 3268 385 3271
rect 662 3271 665 3281
rect 1018 3278 1025 3281
rect 646 3268 665 3271
rect 750 3268 761 3271
rect 950 3268 958 3271
rect 1110 3271 1113 3281
rect 1158 3278 1174 3281
rect 1358 3278 1377 3281
rect 1662 3278 1681 3281
rect 1158 3274 1162 3278
rect 1110 3268 1129 3271
rect 1230 3268 1242 3271
rect 1814 3271 1817 3281
rect 1918 3272 1921 3281
rect 2502 3278 2513 3281
rect 2502 3272 2505 3278
rect 2814 3272 2817 3281
rect 3126 3281 3129 3288
rect 3126 3278 3137 3281
rect 1798 3268 1817 3271
rect 2130 3268 2145 3271
rect 2366 3268 2385 3271
rect 3102 3268 3113 3271
rect 3386 3268 3393 3271
rect 22 3258 34 3261
rect 370 3258 377 3261
rect 758 3262 761 3268
rect 886 3258 889 3268
rect 1006 3261 1009 3268
rect 978 3258 985 3261
rect 990 3258 1009 3261
rect 1134 3258 1146 3261
rect 1574 3258 1590 3261
rect 1782 3258 1790 3261
rect 1862 3258 1881 3261
rect 1894 3258 1913 3261
rect 2078 3261 2081 3268
rect 2070 3258 2081 3261
rect 2562 3258 2569 3261
rect 2698 3258 2705 3261
rect 2822 3258 2830 3261
rect 3110 3262 3113 3268
rect 3374 3258 3382 3261
rect 3502 3258 3510 3261
rect 30 3257 34 3258
rect 1142 3257 1146 3258
rect 1782 3257 1786 3258
rect 1506 3248 1510 3252
rect 1878 3248 1881 3258
rect 1890 3248 1894 3252
rect 562 3238 565 3242
rect 1069 3238 1070 3242
rect 1763 3238 1766 3242
rect 2206 3241 2209 3251
rect 2842 3248 2846 3252
rect 2198 3238 2209 3241
rect 2250 3228 2251 3232
rect 3402 3228 3403 3232
rect 970 3218 971 3222
rect 480 3203 482 3207
rect 486 3203 489 3207
rect 493 3203 496 3207
rect 1512 3203 1514 3207
rect 1518 3203 1521 3207
rect 1525 3203 1528 3207
rect 2536 3203 2538 3207
rect 2542 3203 2545 3207
rect 2549 3203 2552 3207
rect 933 3188 934 3192
rect 1837 3188 1838 3192
rect 3298 3188 3299 3192
rect 70 3168 81 3171
rect 818 3168 819 3172
rect 1205 3168 1206 3172
rect 1398 3168 1406 3171
rect 78 3162 81 3168
rect 62 3151 65 3161
rect 586 3158 590 3162
rect 1314 3158 1316 3162
rect 2286 3158 2297 3161
rect 2498 3158 2505 3161
rect 46 3148 65 3151
rect 246 3148 254 3151
rect 410 3148 425 3151
rect 478 3148 494 3151
rect 510 3148 521 3151
rect 770 3148 785 3151
rect 870 3148 889 3151
rect 934 3148 961 3151
rect 178 3138 193 3141
rect 198 3138 206 3141
rect 405 3138 406 3142
rect 522 3138 529 3141
rect 534 3138 542 3141
rect 606 3138 617 3141
rect 646 3138 654 3141
rect 798 3138 801 3148
rect 1122 3148 1129 3151
rect 1174 3148 1190 3151
rect 1206 3148 1225 3151
rect 1446 3148 1457 3151
rect 1574 3151 1578 3153
rect 2294 3152 2297 3158
rect 3054 3153 3058 3158
rect 1574 3148 1585 3151
rect 1666 3148 1673 3151
rect 1746 3148 1753 3151
rect 1782 3148 1793 3151
rect 1850 3148 1865 3151
rect 1702 3141 1705 3148
rect 1782 3142 1785 3148
rect 1998 3148 2006 3151
rect 2198 3148 2217 3151
rect 2438 3151 2442 3153
rect 1702 3138 1713 3141
rect 1734 3138 1742 3141
rect 2158 3138 2166 3141
rect 2274 3138 2281 3141
rect 2314 3138 2321 3141
rect 2342 3138 2345 3148
rect 2438 3148 2449 3151
rect 2754 3148 2761 3151
rect 2950 3148 2958 3151
rect 3206 3151 3210 3153
rect 3206 3148 3217 3151
rect 3302 3148 3321 3151
rect 2726 3138 2745 3141
rect 2806 3138 2825 3141
rect 3082 3138 3105 3141
rect 3246 3138 3265 3141
rect 3358 3138 3369 3141
rect 3506 3138 3513 3141
rect 3550 3138 3558 3141
rect 334 3128 353 3131
rect 534 3128 537 3138
rect 606 3132 609 3138
rect 646 3128 649 3138
rect 682 3128 689 3131
rect 698 3128 705 3131
rect 758 3128 766 3131
rect 1354 3128 1361 3131
rect 1414 3128 1425 3131
rect 1762 3128 1769 3131
rect 2126 3128 2134 3131
rect 2806 3128 2809 3138
rect 3358 3132 3361 3138
rect 3274 3128 3289 3131
rect 3398 3131 3401 3138
rect 3406 3131 3410 3133
rect 3398 3128 3410 3131
rect 1636 3118 1638 3122
rect 2266 3118 2267 3122
rect 2301 3118 2302 3122
rect 3070 3118 3078 3121
rect 992 3103 994 3107
rect 998 3103 1001 3107
rect 1005 3103 1008 3107
rect 2024 3103 2026 3107
rect 2030 3103 2033 3107
rect 2037 3103 2040 3107
rect 3040 3103 3042 3107
rect 3046 3103 3049 3107
rect 3053 3103 3056 3107
rect 498 3088 505 3091
rect 1461 3088 1462 3092
rect 1956 3088 1958 3092
rect 14 3078 22 3081
rect 78 3071 81 3081
rect 302 3078 321 3081
rect 78 3068 97 3071
rect 102 3068 113 3071
rect 390 3071 393 3081
rect 2030 3078 2046 3081
rect 374 3068 393 3071
rect 406 3068 425 3071
rect 446 3068 457 3071
rect 742 3068 761 3071
rect 806 3068 825 3071
rect 838 3068 857 3071
rect 878 3068 897 3071
rect 1154 3068 1169 3071
rect 1182 3068 1201 3071
rect 1318 3068 1326 3071
rect 1586 3068 1601 3071
rect 1750 3068 1758 3071
rect 1850 3068 1857 3071
rect 1890 3068 1897 3071
rect 2054 3071 2057 3081
rect 2018 3068 2057 3071
rect 2206 3068 2225 3071
rect 2278 3068 2289 3071
rect 2398 3068 2409 3071
rect 2846 3071 2849 3081
rect 2966 3078 2974 3081
rect 3066 3078 3081 3081
rect 2966 3077 2970 3078
rect 2846 3068 2865 3071
rect 3370 3068 3377 3071
rect 102 3062 105 3068
rect 454 3062 457 3068
rect 262 3058 281 3061
rect 838 3062 841 3068
rect 962 3058 977 3061
rect 1250 3058 1265 3061
rect 1314 3058 1337 3061
rect 1534 3058 1553 3061
rect 1574 3058 1593 3061
rect 1702 3061 1705 3068
rect 1686 3058 1705 3061
rect 1730 3058 1737 3061
rect 1862 3058 1873 3061
rect 1910 3058 1926 3061
rect 2174 3058 2185 3061
rect 2270 3061 2273 3068
rect 2254 3058 2273 3061
rect 2286 3062 2289 3068
rect 2406 3062 2409 3068
rect 2458 3058 2465 3061
rect 2966 3058 2977 3061
rect 3070 3061 3073 3068
rect 3046 3058 3073 3061
rect 3214 3058 3217 3068
rect 3326 3058 3345 3061
rect 3350 3058 3369 3061
rect 3430 3058 3438 3061
rect 3486 3058 3497 3061
rect 2966 3057 2970 3058
rect 3486 3057 3490 3058
rect 166 3048 185 3051
rect 638 3048 657 3051
rect 794 3048 798 3052
rect 990 3048 1017 3051
rect 2234 3048 2241 3051
rect 710 3038 718 3041
rect 949 3038 950 3042
rect 1309 3038 1310 3042
rect 1381 3028 1382 3032
rect 669 3018 670 3022
rect 746 3018 747 3022
rect 978 3018 979 3022
rect 1362 3018 1363 3022
rect 2253 3018 2254 3022
rect 2981 3018 2982 3022
rect 480 3003 482 3007
rect 486 3003 489 3007
rect 493 3003 496 3007
rect 1512 3003 1514 3007
rect 1518 3003 1521 3007
rect 1525 3003 1528 3007
rect 2536 3003 2538 3007
rect 2542 3003 2545 3007
rect 2549 3003 2552 3007
rect 173 2988 174 2992
rect 285 2988 286 2992
rect 354 2988 355 2992
rect 466 2988 467 2992
rect 522 2988 523 2992
rect 1117 2988 1118 2992
rect 2106 2988 2107 2992
rect 2530 2988 2531 2992
rect 2845 2988 2846 2992
rect 2954 2988 2955 2992
rect 2986 2988 2987 2992
rect 3226 2988 3227 2992
rect 1349 2978 1350 2982
rect 534 2968 545 2971
rect 890 2968 897 2971
rect 1294 2968 1302 2971
rect 2562 2968 2569 2971
rect 1366 2958 1385 2961
rect 1390 2958 1409 2961
rect 1486 2958 1505 2961
rect 1530 2958 1545 2961
rect 1930 2958 1937 2961
rect 2170 2958 2174 2962
rect 2330 2958 2337 2961
rect 30 2948 49 2951
rect 22 2938 38 2941
rect 166 2941 169 2951
rect 286 2948 305 2951
rect 314 2948 321 2951
rect 422 2948 438 2951
rect 486 2948 521 2951
rect 562 2948 569 2951
rect 150 2938 169 2941
rect 186 2938 201 2941
rect 222 2938 241 2941
rect 406 2941 409 2948
rect 622 2942 625 2951
rect 654 2948 665 2951
rect 806 2948 833 2951
rect 1070 2948 1078 2951
rect 1122 2948 1145 2951
rect 1270 2948 1297 2951
rect 1478 2948 1489 2951
rect 1562 2948 1577 2951
rect 1758 2948 1766 2951
rect 2046 2948 2054 2951
rect 2302 2951 2305 2958
rect 2430 2951 2434 2953
rect 2294 2948 2305 2951
rect 406 2938 417 2941
rect 506 2938 513 2941
rect 610 2938 617 2941
rect 842 2938 857 2941
rect 934 2938 950 2941
rect 1074 2938 1089 2941
rect 1254 2938 1257 2948
rect 1518 2938 1534 2941
rect 1574 2938 1577 2948
rect 1894 2938 1897 2948
rect 2430 2948 2441 2951
rect 2458 2948 2473 2951
rect 2510 2948 2518 2951
rect 2610 2948 2625 2951
rect 2678 2948 2686 2951
rect 2702 2948 2710 2951
rect 2998 2951 3001 2961
rect 2998 2948 3017 2951
rect 3314 2948 3321 2951
rect 1962 2938 1969 2941
rect 1974 2938 1982 2941
rect 2010 2938 2038 2941
rect 2262 2938 2289 2941
rect 2894 2938 2918 2941
rect 3078 2938 3086 2941
rect 3110 2938 3126 2941
rect 3162 2938 3169 2941
rect 3326 2941 3329 2951
rect 3342 2948 3361 2951
rect 3414 2948 3430 2951
rect 3542 2948 3550 2951
rect 3326 2938 3345 2941
rect 170 2928 177 2931
rect 182 2928 190 2931
rect 310 2928 329 2931
rect 558 2928 566 2931
rect 834 2928 838 2932
rect 910 2928 918 2931
rect 1694 2928 1713 2931
rect 2438 2931 2441 2938
rect 2438 2928 2449 2931
rect 3482 2928 3489 2931
rect 3494 2928 3502 2931
rect 3522 2928 3529 2931
rect 858 2918 859 2922
rect 1660 2918 1662 2922
rect 2229 2918 2230 2922
rect 2309 2918 2310 2922
rect 3054 2921 3057 2928
rect 3046 2918 3057 2921
rect 992 2903 994 2907
rect 998 2903 1001 2907
rect 1005 2903 1008 2907
rect 2024 2903 2026 2907
rect 2030 2903 2033 2907
rect 2037 2903 2040 2907
rect 3040 2903 3042 2907
rect 3046 2903 3049 2907
rect 3053 2903 3056 2907
rect 1221 2888 1222 2892
rect 1338 2888 1339 2892
rect 2373 2888 2374 2892
rect 26 2878 33 2881
rect 62 2878 70 2881
rect 102 2878 110 2881
rect 438 2878 446 2881
rect 714 2878 726 2881
rect 778 2878 785 2881
rect 818 2878 825 2881
rect 1030 2872 1033 2881
rect 1262 2878 1270 2881
rect 1482 2878 1486 2882
rect 1958 2878 1969 2881
rect 2114 2878 2121 2882
rect 1966 2872 1969 2878
rect 2118 2872 2121 2878
rect 2638 2872 2641 2881
rect 2962 2878 2978 2881
rect 3010 2878 3017 2882
rect 3198 2878 3209 2881
rect 2974 2874 2978 2878
rect 3014 2872 3017 2878
rect 3206 2872 3209 2878
rect 174 2868 185 2871
rect 222 2868 230 2871
rect 246 2868 257 2871
rect 330 2868 337 2871
rect 386 2868 393 2871
rect 174 2862 177 2868
rect 22 2858 49 2861
rect 246 2858 254 2861
rect 326 2858 334 2861
rect 462 2858 478 2861
rect 518 2861 521 2871
rect 702 2868 718 2871
rect 758 2868 785 2871
rect 1094 2868 1102 2871
rect 1166 2868 1174 2871
rect 1398 2868 1406 2871
rect 1434 2868 1441 2871
rect 1498 2868 1521 2871
rect 1662 2868 1681 2871
rect 1850 2868 1865 2871
rect 2142 2868 2158 2871
rect 518 2858 529 2861
rect 606 2858 633 2861
rect 938 2858 953 2861
rect 958 2858 977 2861
rect 1002 2858 1009 2861
rect 1062 2858 1070 2861
rect 1166 2858 1169 2868
rect 1178 2858 1185 2861
rect 1438 2858 1441 2868
rect 2018 2858 2033 2861
rect 2062 2858 2070 2861
rect 2102 2861 2105 2868
rect 2086 2858 2105 2861
rect 2174 2858 2185 2861
rect 2246 2858 2265 2861
rect 2270 2858 2278 2861
rect 2290 2858 2297 2861
rect 2342 2861 2345 2871
rect 2506 2868 2513 2871
rect 2538 2868 2553 2871
rect 3290 2868 3305 2871
rect 3322 2868 3329 2871
rect 3390 2871 3393 2881
rect 3362 2868 3369 2871
rect 3374 2868 3393 2871
rect 3462 2868 3470 2871
rect 3518 2868 3526 2871
rect 2334 2858 2345 2861
rect 2350 2858 2358 2861
rect 2798 2858 2806 2861
rect 3110 2858 3137 2861
rect 3142 2858 3161 2861
rect 3174 2858 3190 2861
rect 3266 2858 3281 2861
rect 202 2848 209 2851
rect 409 2848 414 2852
rect 1230 2851 1233 2858
rect 1230 2848 1241 2851
rect 1286 2848 1297 2851
rect 1612 2848 1614 2852
rect 1930 2848 1937 2851
rect 2118 2851 2121 2858
rect 2174 2852 2177 2858
rect 2334 2856 2338 2858
rect 2118 2848 2129 2851
rect 3158 2848 3161 2858
rect 670 2841 673 2848
rect 2806 2842 2810 2844
rect 662 2838 673 2841
rect 1746 2838 1753 2841
rect 3022 2838 3054 2841
rect 925 2828 926 2832
rect 133 2818 134 2822
rect 373 2818 374 2822
rect 509 2818 510 2822
rect 637 2818 638 2822
rect 853 2818 854 2822
rect 893 2818 894 2822
rect 1133 2818 1134 2822
rect 1805 2818 1806 2822
rect 1997 2818 1998 2822
rect 2085 2818 2086 2822
rect 2189 2818 2190 2822
rect 2589 2818 2590 2822
rect 2829 2818 2830 2822
rect 3093 2818 3094 2822
rect 3173 2818 3174 2822
rect 480 2803 482 2807
rect 486 2803 489 2807
rect 493 2803 496 2807
rect 1512 2803 1514 2807
rect 1518 2803 1521 2807
rect 1525 2803 1528 2807
rect 2536 2803 2538 2807
rect 2542 2803 2545 2807
rect 2549 2803 2552 2807
rect 34 2788 35 2792
rect 117 2788 118 2792
rect 2006 2788 2022 2791
rect 2301 2788 2302 2792
rect 2485 2788 2486 2792
rect 2565 2788 2566 2792
rect 2794 2788 2795 2792
rect 246 2768 258 2771
rect 954 2768 969 2771
rect 1798 2768 1809 2771
rect 2109 2768 2110 2772
rect 3474 2768 3475 2772
rect 1806 2762 1809 2768
rect 94 2758 105 2761
rect 266 2758 270 2762
rect 382 2758 393 2761
rect 518 2758 537 2761
rect 1538 2758 1545 2761
rect 118 2748 142 2751
rect 162 2748 169 2751
rect 202 2748 209 2751
rect 282 2748 289 2751
rect 354 2748 369 2751
rect 374 2748 382 2751
rect 446 2748 454 2751
rect 498 2748 505 2751
rect 574 2748 585 2751
rect 646 2748 657 2751
rect 806 2748 814 2751
rect 1174 2748 1182 2751
rect 1294 2751 1298 2753
rect 582 2742 585 2748
rect 1294 2748 1305 2751
rect 1510 2748 1545 2751
rect 1614 2751 1617 2761
rect 1670 2758 1689 2761
rect 1742 2758 1753 2761
rect 1942 2758 1953 2761
rect 1962 2758 1966 2762
rect 2086 2758 2097 2761
rect 1598 2748 1617 2751
rect 1662 2748 1673 2751
rect 1766 2748 1782 2751
rect 1978 2748 1985 2751
rect 2134 2748 2153 2751
rect 2206 2748 2222 2751
rect 2522 2748 2550 2751
rect 2658 2748 2670 2751
rect 2830 2751 2833 2761
rect 2870 2758 2881 2761
rect 2830 2748 2841 2751
rect 3118 2748 3134 2751
rect 3270 2748 3278 2751
rect 3426 2748 3441 2751
rect 3478 2748 3486 2751
rect 2838 2742 2841 2748
rect 126 2738 134 2741
rect 174 2738 182 2741
rect 206 2738 217 2741
rect 330 2738 345 2741
rect 442 2738 465 2741
rect 734 2738 753 2741
rect 810 2738 817 2741
rect 878 2738 886 2741
rect 902 2738 910 2741
rect 972 2738 974 2742
rect 1302 2738 1313 2741
rect 1558 2738 1569 2741
rect 1898 2738 1905 2741
rect 2310 2738 2321 2741
rect 2590 2738 2609 2741
rect 2622 2738 2649 2741
rect 2686 2738 2697 2741
rect 2790 2738 2801 2741
rect 2910 2738 2918 2741
rect 3226 2738 3249 2741
rect 78 2728 89 2731
rect 174 2728 177 2738
rect 206 2732 209 2738
rect 1302 2732 1305 2738
rect 1566 2732 1569 2738
rect 586 2728 593 2731
rect 1038 2728 1049 2731
rect 1886 2728 1897 2731
rect 2606 2728 2609 2738
rect 2798 2732 2801 2738
rect 3058 2728 3065 2731
rect 194 2718 195 2722
rect 1122 2718 1123 2722
rect 1818 2718 1819 2722
rect 2724 2718 2726 2722
rect 992 2703 994 2707
rect 998 2703 1001 2707
rect 1005 2703 1008 2707
rect 2024 2703 2026 2707
rect 2030 2703 2033 2707
rect 2037 2703 2040 2707
rect 3040 2703 3042 2707
rect 3046 2703 3049 2707
rect 3053 2703 3056 2707
rect 434 2688 435 2692
rect 1045 2688 1046 2692
rect 2477 2688 2478 2692
rect 2674 2688 2675 2692
rect 3050 2688 3057 2691
rect 3306 2688 3308 2692
rect 3316 2688 3318 2692
rect 54 2668 62 2671
rect 78 2671 81 2678
rect 70 2668 81 2671
rect 290 2668 305 2671
rect 358 2671 361 2681
rect 778 2678 793 2681
rect 1734 2678 1753 2681
rect 2554 2678 2561 2681
rect 2910 2678 2918 2682
rect 342 2668 361 2671
rect 366 2668 390 2671
rect 454 2668 473 2671
rect 822 2668 841 2671
rect 954 2668 969 2671
rect 1198 2668 1209 2671
rect 10 2658 17 2661
rect 86 2658 94 2661
rect 122 2658 137 2661
rect 246 2658 262 2661
rect 758 2661 761 2668
rect 750 2658 761 2661
rect 790 2658 798 2661
rect 946 2658 961 2661
rect 982 2658 1009 2661
rect 1110 2658 1113 2668
rect 1206 2662 1209 2668
rect 1438 2668 1454 2671
rect 1502 2668 1510 2671
rect 1546 2668 1553 2671
rect 1618 2668 1633 2671
rect 1698 2668 1705 2671
rect 1910 2668 1921 2671
rect 1950 2668 1961 2671
rect 2114 2668 2121 2671
rect 2162 2668 2169 2671
rect 2206 2668 2214 2671
rect 2350 2668 2369 2671
rect 1918 2662 1921 2668
rect 1242 2658 1249 2661
rect 1862 2658 1889 2661
rect 1998 2658 2006 2661
rect 2078 2658 2089 2661
rect 2174 2658 2193 2661
rect 2270 2658 2289 2661
rect 2294 2658 2302 2661
rect 2374 2658 2393 2661
rect 2398 2658 2401 2678
rect 2454 2668 2470 2671
rect 2486 2661 2489 2671
rect 2534 2668 2558 2671
rect 2846 2671 2849 2678
rect 2910 2672 2913 2678
rect 2846 2668 2857 2671
rect 3022 2668 3030 2671
rect 3078 2668 3089 2671
rect 3110 2668 3118 2671
rect 2486 2658 2494 2661
rect 2514 2658 2521 2661
rect 2538 2658 2569 2661
rect 2670 2658 2689 2661
rect 2702 2658 2729 2661
rect 2902 2658 2910 2661
rect 2930 2658 2937 2661
rect 3134 2661 3137 2668
rect 3126 2658 3137 2661
rect 3202 2658 3217 2661
rect 3250 2658 3257 2661
rect 1462 2648 1481 2651
rect 2038 2648 2049 2651
rect 2502 2648 2513 2651
rect 2686 2648 2689 2658
rect 3126 2648 3137 2651
rect 3470 2648 3481 2651
rect 706 2638 707 2642
rect 814 2638 822 2641
rect 1122 2638 1134 2641
rect 2038 2641 2041 2648
rect 2022 2638 2041 2641
rect 3514 2638 3516 2642
rect 906 2628 907 2632
rect 138 2618 139 2622
rect 570 2618 571 2622
rect 858 2618 859 2622
rect 1493 2618 1494 2622
rect 1562 2618 1563 2622
rect 2266 2618 2267 2622
rect 2314 2618 2315 2622
rect 2341 2618 2342 2622
rect 480 2603 482 2607
rect 486 2603 489 2607
rect 493 2603 496 2607
rect 1512 2603 1514 2607
rect 1518 2603 1521 2607
rect 1525 2603 1528 2607
rect 2536 2603 2538 2607
rect 2542 2603 2545 2607
rect 2549 2603 2552 2607
rect 101 2588 102 2592
rect 226 2588 227 2592
rect 261 2588 262 2592
rect 597 2588 598 2592
rect 685 2588 686 2592
rect 749 2588 750 2592
rect 1842 2588 1843 2592
rect 1973 2588 1974 2592
rect 2429 2588 2430 2592
rect 2717 2588 2718 2592
rect 3285 2588 3286 2592
rect 3404 2588 3406 2592
rect 2581 2578 2582 2582
rect 3542 2578 3550 2581
rect 1070 2568 1078 2571
rect 2813 2568 2814 2572
rect 2962 2568 2963 2572
rect 3058 2568 3065 2571
rect 3354 2568 3361 2571
rect 782 2566 786 2568
rect 1070 2566 1074 2568
rect 1278 2566 1282 2568
rect 86 2548 97 2551
rect 114 2548 121 2551
rect 138 2548 145 2551
rect 238 2551 241 2561
rect 654 2558 665 2561
rect 862 2558 870 2561
rect 2198 2558 2217 2561
rect 2318 2558 2329 2561
rect 238 2548 257 2551
rect 566 2551 569 2558
rect 2486 2552 2489 2561
rect 2694 2558 2705 2561
rect 558 2548 569 2551
rect 662 2548 681 2551
rect 750 2548 766 2551
rect 794 2548 801 2551
rect 1146 2548 1153 2551
rect 1190 2548 1209 2551
rect 162 2538 169 2541
rect 374 2541 377 2548
rect 366 2538 377 2541
rect 630 2538 641 2541
rect 1126 2538 1134 2541
rect 1174 2541 1177 2548
rect 1166 2538 1177 2541
rect 1430 2541 1433 2551
rect 1974 2548 2001 2551
rect 2042 2548 2057 2551
rect 2118 2548 2137 2551
rect 2190 2548 2201 2551
rect 2218 2548 2225 2551
rect 2230 2548 2249 2551
rect 2290 2548 2305 2551
rect 2430 2548 2457 2551
rect 2522 2548 2529 2551
rect 2798 2551 2801 2561
rect 2718 2548 2745 2551
rect 2766 2548 2777 2551
rect 2782 2548 2801 2551
rect 2814 2548 2833 2551
rect 2974 2551 2977 2561
rect 2974 2548 2993 2551
rect 3322 2548 3329 2551
rect 3462 2548 3470 2551
rect 3518 2551 3522 2553
rect 3518 2548 3529 2551
rect 1430 2538 1438 2541
rect 1502 2538 1526 2541
rect 1534 2538 1542 2541
rect 1750 2538 1766 2541
rect 2022 2538 2038 2541
rect 2190 2542 2193 2548
rect 2142 2538 2150 2541
rect 2490 2538 2497 2541
rect 2518 2538 2521 2548
rect 2650 2538 2657 2541
rect 3086 2538 3094 2541
rect 3174 2538 3193 2541
rect 3310 2538 3321 2541
rect 630 2532 633 2538
rect 86 2528 94 2531
rect 414 2528 433 2531
rect 1422 2528 1430 2531
rect 1522 2528 1529 2531
rect 2014 2531 2017 2538
rect 2002 2528 2017 2531
rect 2034 2528 2046 2531
rect 2142 2528 2145 2538
rect 2526 2531 2529 2538
rect 2526 2528 2537 2531
rect 2910 2528 2921 2531
rect 3174 2528 3177 2538
rect 3310 2532 3313 2538
rect 3218 2528 3230 2531
rect 3294 2528 3305 2531
rect 578 2518 579 2522
rect 778 2518 779 2522
rect 858 2518 859 2522
rect 909 2518 910 2522
rect 1066 2518 1067 2522
rect 1274 2518 1275 2522
rect 1493 2518 1494 2522
rect 1773 2518 1774 2522
rect 992 2503 994 2507
rect 998 2503 1001 2507
rect 1005 2503 1008 2507
rect 2024 2503 2026 2507
rect 2030 2503 2033 2507
rect 2037 2503 2040 2507
rect 3040 2503 3042 2507
rect 3046 2503 3049 2507
rect 3053 2503 3056 2507
rect 2301 2488 2302 2492
rect 3474 2488 3475 2492
rect 702 2478 713 2481
rect 1798 2478 1806 2481
rect 98 2468 105 2471
rect 318 2468 337 2471
rect 366 2468 374 2471
rect 654 2468 662 2471
rect 734 2468 742 2471
rect 30 2458 38 2461
rect 86 2458 102 2461
rect 370 2458 385 2461
rect 486 2458 510 2461
rect 558 2458 574 2461
rect 590 2458 598 2461
rect 646 2458 670 2461
rect 862 2458 870 2461
rect 1010 2458 1033 2461
rect 1070 2461 1073 2471
rect 1066 2458 1073 2461
rect 1078 2458 1097 2461
rect 1110 2458 1118 2461
rect 1214 2458 1233 2461
rect 1278 2458 1286 2461
rect 1342 2461 1345 2471
rect 1318 2458 1337 2461
rect 1342 2458 1358 2461
rect 1478 2458 1486 2461
rect 1558 2461 1561 2471
rect 1606 2468 1614 2471
rect 1690 2468 1697 2471
rect 1710 2468 1729 2471
rect 1870 2468 1889 2471
rect 1946 2468 1953 2471
rect 2006 2468 2014 2471
rect 2134 2468 2145 2471
rect 2462 2471 2465 2481
rect 2638 2478 2657 2481
rect 3198 2478 3209 2481
rect 2446 2468 2465 2471
rect 2486 2468 2505 2471
rect 2562 2468 2577 2471
rect 1558 2458 1574 2461
rect 1802 2458 1809 2461
rect 1886 2458 1889 2468
rect 2134 2462 2137 2468
rect 2014 2458 2041 2461
rect 2486 2458 2489 2468
rect 2554 2458 2569 2461
rect 2614 2458 2630 2461
rect 2634 2458 2641 2461
rect 2658 2458 2665 2461
rect 2710 2461 2713 2471
rect 2756 2468 2758 2472
rect 2858 2468 2865 2471
rect 2958 2468 2969 2471
rect 2982 2468 3001 2471
rect 3438 2471 3441 2481
rect 3402 2468 3417 2471
rect 3422 2468 3441 2471
rect 3446 2468 3465 2471
rect 3486 2468 3505 2471
rect 2966 2462 2969 2468
rect 2698 2458 2713 2461
rect 2718 2458 2726 2461
rect 2770 2458 2777 2461
rect 3006 2458 3014 2461
rect 3094 2458 3102 2461
rect 3110 2458 3121 2461
rect 3270 2458 3289 2461
rect 3306 2458 3318 2461
rect 3390 2458 3406 2461
rect 3462 2458 3465 2468
rect 3510 2461 3513 2468
rect 3502 2458 3513 2461
rect 30 2448 33 2458
rect 121 2448 126 2452
rect 246 2448 265 2451
rect 502 2448 529 2451
rect 614 2448 633 2451
rect 766 2451 769 2458
rect 766 2448 785 2451
rect 1094 2448 1097 2458
rect 1230 2448 1233 2458
rect 1318 2448 1321 2458
rect 1518 2448 1526 2451
rect 2982 2451 2985 2458
rect 3118 2452 3121 2458
rect 2974 2448 2985 2451
rect 3026 2448 3030 2452
rect 3286 2448 3289 2458
rect 502 2442 505 2448
rect 2750 2446 2754 2448
rect 454 2438 462 2441
rect 1486 2438 1510 2441
rect 1550 2438 1558 2441
rect 1765 2438 1766 2442
rect 2542 2438 2550 2441
rect 2738 2438 2753 2441
rect 1141 2428 1142 2432
rect 18 2418 19 2422
rect 397 2418 398 2422
rect 437 2418 438 2422
rect 485 2418 486 2422
rect 557 2418 558 2422
rect 645 2418 646 2422
rect 674 2418 675 2422
rect 754 2418 755 2422
rect 821 2418 822 2422
rect 861 2418 862 2422
rect 1045 2418 1046 2422
rect 1109 2418 1110 2422
rect 1181 2418 1182 2422
rect 1245 2418 1246 2422
rect 1277 2418 1278 2422
rect 1373 2418 1374 2422
rect 1893 2418 1894 2422
rect 1925 2418 1926 2422
rect 3250 2418 3251 2422
rect 480 2403 482 2407
rect 486 2403 489 2407
rect 493 2403 496 2407
rect 1512 2403 1514 2407
rect 1518 2403 1521 2407
rect 1525 2403 1528 2407
rect 2536 2403 2538 2407
rect 2542 2403 2545 2407
rect 2549 2403 2552 2407
rect 2405 2388 2406 2392
rect 2738 2388 2739 2392
rect 3093 2388 3094 2392
rect 3394 2388 3395 2392
rect 346 2368 347 2372
rect 606 2368 614 2371
rect 734 2368 745 2371
rect 2234 2368 2235 2372
rect 2290 2368 2297 2371
rect 2788 2368 2790 2372
rect 2938 2368 2939 2372
rect 3292 2368 3294 2372
rect 406 2366 410 2368
rect 734 2362 737 2368
rect 326 2351 329 2361
rect 438 2358 457 2361
rect 486 2358 502 2361
rect 990 2358 998 2361
rect 326 2348 342 2351
rect 410 2348 425 2351
rect 638 2351 641 2358
rect 622 2348 641 2351
rect 674 2348 681 2351
rect 794 2348 801 2351
rect 878 2348 886 2351
rect 982 2348 998 2351
rect 1062 2351 1065 2361
rect 1062 2348 1081 2351
rect 1182 2348 1190 2351
rect 1222 2351 1225 2361
rect 1206 2348 1225 2351
rect 1250 2348 1265 2351
rect 1382 2351 1385 2361
rect 1518 2358 1529 2361
rect 1590 2358 1598 2361
rect 1614 2358 1625 2361
rect 1366 2348 1385 2351
rect 1454 2351 1457 2358
rect 1526 2352 1529 2358
rect 1614 2352 1617 2358
rect 1446 2348 1457 2351
rect 1478 2348 1497 2351
rect 1538 2348 1545 2351
rect 1622 2348 1641 2351
rect 1646 2348 1657 2351
rect 1710 2351 1713 2361
rect 1974 2358 1982 2361
rect 2078 2358 2089 2361
rect 2158 2361 2161 2368
rect 2158 2358 2169 2361
rect 3074 2358 3081 2361
rect 3178 2358 3185 2361
rect 1710 2348 1729 2351
rect 1934 2348 1961 2351
rect 1974 2348 1993 2351
rect 2010 2348 2017 2351
rect 2022 2348 2038 2351
rect 2134 2348 2153 2351
rect 2190 2348 2198 2351
rect 2278 2351 2282 2354
rect 2262 2348 2282 2351
rect 2310 2348 2318 2351
rect 2406 2348 2414 2351
rect 2474 2348 2489 2351
rect 2614 2348 2622 2351
rect 2722 2348 2734 2351
rect 2834 2348 2849 2351
rect 202 2338 209 2341
rect 262 2338 273 2341
rect 306 2338 313 2341
rect 574 2338 582 2341
rect 822 2338 825 2348
rect 878 2338 881 2348
rect 1654 2342 1657 2348
rect 1194 2338 1201 2341
rect 1246 2338 1254 2341
rect 1306 2338 1313 2341
rect 1606 2338 1614 2341
rect 1670 2338 1689 2341
rect 1782 2341 1785 2348
rect 1782 2338 1793 2341
rect 1866 2338 1873 2341
rect 2322 2338 2329 2341
rect 2526 2338 2569 2341
rect 2614 2338 2617 2348
rect 2846 2338 2849 2348
rect 2894 2341 2897 2351
rect 2962 2348 2969 2351
rect 3030 2348 3041 2351
rect 3150 2348 3158 2351
rect 3186 2348 3193 2351
rect 3198 2348 3214 2351
rect 3386 2348 3393 2351
rect 3530 2348 3537 2351
rect 3038 2342 3041 2348
rect 2894 2338 2913 2341
rect 2974 2338 2993 2341
rect 3002 2338 3017 2341
rect 3162 2338 3169 2341
rect 3210 2338 3217 2341
rect 3442 2338 3449 2341
rect 3470 2338 3489 2341
rect 3502 2338 3521 2341
rect 3550 2338 3558 2341
rect 1902 2328 1910 2331
rect 1958 2328 1966 2331
rect 2110 2328 2113 2338
rect 2134 2331 2137 2338
rect 2134 2328 2150 2331
rect 2666 2328 2670 2332
rect 2998 2328 3006 2331
rect 293 2318 294 2322
rect 373 2318 374 2322
rect 402 2318 403 2322
rect 538 2318 539 2322
rect 2205 2318 2206 2322
rect 2300 2318 2302 2322
rect 2452 2318 2454 2322
rect 992 2303 994 2307
rect 998 2303 1001 2307
rect 1005 2303 1008 2307
rect 2024 2303 2026 2307
rect 2030 2303 2033 2307
rect 2037 2303 2040 2307
rect 3040 2303 3042 2307
rect 3046 2303 3049 2307
rect 3053 2303 3056 2307
rect 50 2288 51 2292
rect 2117 2288 2118 2292
rect 2550 2288 2566 2291
rect 2645 2288 2646 2292
rect 2781 2288 2782 2292
rect 3314 2288 3315 2292
rect 3333 2288 3334 2292
rect 22 2258 30 2261
rect 46 2258 65 2261
rect 78 2258 94 2261
rect 234 2258 241 2261
rect 282 2258 289 2261
rect 318 2261 321 2271
rect 362 2268 369 2271
rect 306 2258 321 2261
rect 430 2261 433 2281
rect 574 2272 577 2281
rect 1498 2278 1505 2281
rect 1738 2278 1745 2282
rect 1974 2278 1982 2281
rect 2174 2278 2185 2281
rect 2202 2278 2209 2281
rect 2814 2278 2825 2281
rect 430 2258 438 2261
rect 454 2258 462 2261
rect 718 2258 737 2261
rect 870 2258 889 2261
rect 1018 2258 1041 2261
rect 1086 2261 1089 2271
rect 1174 2268 1182 2271
rect 1470 2271 1473 2278
rect 1742 2272 1745 2278
rect 1462 2268 1473 2271
rect 1694 2268 1702 2271
rect 1846 2271 1849 2278
rect 2182 2272 2185 2278
rect 2814 2272 2817 2278
rect 1846 2268 1865 2271
rect 1982 2268 1998 2271
rect 2214 2268 2230 2271
rect 1086 2258 1094 2261
rect 1098 2258 1105 2261
rect 1134 2258 1142 2261
rect 1178 2258 1193 2261
rect 1298 2258 1313 2261
rect 1358 2258 1377 2261
rect 1470 2258 1478 2261
rect 1486 2258 1497 2261
rect 1638 2258 1646 2261
rect 1654 2258 1673 2261
rect 1686 2258 1713 2261
rect 1742 2258 1761 2261
rect 1982 2258 1985 2268
rect 2290 2268 2297 2271
rect 2326 2268 2353 2271
rect 2442 2268 2449 2271
rect 2622 2268 2630 2271
rect 2654 2268 2673 2271
rect 2790 2268 2809 2271
rect 2094 2258 2121 2261
rect 2714 2258 2729 2261
rect 2738 2258 2753 2261
rect 2878 2258 2897 2261
rect 3002 2258 3017 2261
rect 3078 2258 3097 2261
rect 3110 2261 3113 2271
rect 3266 2268 3273 2271
rect 3294 2268 3302 2271
rect 3358 2268 3369 2271
rect 3454 2262 3457 2271
rect 3110 2258 3129 2261
rect 3218 2258 3225 2261
rect 3254 2258 3273 2261
rect 3310 2258 3329 2261
rect 3514 2258 3521 2261
rect 62 2248 65 2258
rect 286 2248 289 2258
rect 434 2248 441 2251
rect 702 2248 721 2251
rect 734 2248 737 2258
rect 886 2248 889 2258
rect 1374 2248 1377 2258
rect 1670 2248 1673 2258
rect 1742 2252 1745 2258
rect 2246 2248 2257 2251
rect 2878 2248 2881 2258
rect 3066 2248 3070 2252
rect 3078 2248 3081 2258
rect 3134 2251 3137 2258
rect 3126 2248 3137 2251
rect 3270 2248 3273 2258
rect 3326 2248 3329 2258
rect 3406 2248 3417 2251
rect 3434 2248 3441 2251
rect 3446 2248 3454 2251
rect 54 2242 58 2244
rect 590 2241 593 2248
rect 726 2242 730 2244
rect 2254 2242 2257 2248
rect 590 2238 601 2241
rect 662 2238 670 2241
rect 690 2238 691 2242
rect 1940 2238 1942 2242
rect 2198 2238 2206 2241
rect 3226 2238 3227 2242
rect 21 2218 22 2222
rect 77 2218 78 2222
rect 165 2218 166 2222
rect 549 2218 550 2222
rect 634 2218 635 2222
rect 749 2218 750 2222
rect 837 2218 838 2222
rect 989 2218 990 2222
rect 1165 2218 1166 2222
rect 1194 2218 1195 2222
rect 1229 2218 1230 2222
rect 1282 2218 1283 2222
rect 1325 2218 1326 2222
rect 1762 2218 1763 2222
rect 2550 2218 2558 2221
rect 2866 2218 2867 2222
rect 2970 2218 2972 2222
rect 3194 2218 3195 2222
rect 480 2203 482 2207
rect 486 2203 489 2207
rect 493 2203 496 2207
rect 1512 2203 1514 2207
rect 1518 2203 1521 2207
rect 1525 2203 1528 2207
rect 2536 2203 2538 2207
rect 2542 2203 2545 2207
rect 2549 2203 2552 2207
rect 1898 2188 1899 2192
rect 1970 2188 1971 2192
rect 2050 2188 2057 2191
rect 2274 2188 2275 2192
rect 3274 2188 3275 2192
rect 3394 2188 3395 2192
rect 1522 2178 1529 2181
rect 3106 2178 3108 2182
rect 2125 2168 2126 2172
rect 2149 2168 2150 2172
rect 410 2158 417 2161
rect 10 2148 17 2151
rect 78 2148 86 2151
rect 150 2151 153 2158
rect 134 2148 153 2151
rect 294 2148 302 2151
rect 394 2148 401 2151
rect 438 2148 454 2151
rect 470 2151 473 2161
rect 534 2158 542 2161
rect 670 2158 678 2161
rect 750 2158 769 2161
rect 778 2158 785 2161
rect 846 2158 854 2161
rect 898 2158 905 2161
rect 990 2158 1025 2161
rect 470 2148 489 2151
rect 718 2151 721 2158
rect 718 2148 737 2151
rect 1054 2151 1057 2158
rect 1142 2151 1145 2161
rect 1038 2148 1057 2151
rect 1126 2148 1145 2151
rect 1226 2148 1241 2151
rect 1374 2151 1377 2158
rect 1406 2151 1409 2161
rect 1926 2158 1937 2161
rect 2818 2158 2822 2162
rect 2930 2158 2934 2162
rect 2950 2158 2958 2161
rect 1290 2148 1297 2151
rect 1374 2148 1393 2151
rect 1406 2148 1425 2151
rect 1494 2148 1518 2151
rect 1606 2151 1609 2158
rect 1590 2148 1609 2151
rect 1702 2151 1706 2152
rect 1686 2148 1706 2151
rect 1914 2148 1929 2151
rect 142 2138 150 2141
rect 302 2138 310 2141
rect 382 2138 390 2141
rect 438 2138 441 2148
rect 494 2138 518 2141
rect 558 2138 566 2141
rect 930 2138 937 2141
rect 1166 2138 1169 2148
rect 1214 2138 1222 2141
rect 1226 2138 1233 2141
rect 1662 2138 1670 2141
rect 1686 2138 1689 2148
rect 2010 2138 2017 2141
rect 2078 2141 2081 2151
rect 2370 2148 2385 2151
rect 2398 2148 2414 2151
rect 2434 2148 2441 2151
rect 2542 2148 2558 2151
rect 2590 2148 2598 2151
rect 2734 2148 2742 2151
rect 2874 2148 2881 2151
rect 2902 2148 2918 2151
rect 2982 2151 2985 2161
rect 3054 2151 3057 2161
rect 3066 2158 3070 2162
rect 2946 2148 2953 2151
rect 2982 2148 3001 2151
rect 3022 2148 3057 2151
rect 3258 2148 3273 2151
rect 3318 2148 3337 2151
rect 3446 2148 3457 2151
rect 2078 2138 2097 2141
rect 2134 2138 2153 2141
rect 2158 2138 2166 2141
rect 2270 2138 2297 2141
rect 2382 2138 2385 2148
rect 2446 2138 2473 2141
rect 2698 2138 2713 2141
rect 3006 2138 3025 2141
rect 346 2128 350 2132
rect 1502 2128 1510 2131
rect 2014 2128 2017 2138
rect 2022 2128 2057 2131
rect 2158 2128 2161 2138
rect 2422 2128 2430 2131
rect 210 2118 211 2122
rect 266 2118 267 2122
rect 666 2118 667 2122
rect 842 2118 843 2122
rect 890 2118 891 2122
rect 909 2118 910 2122
rect 1018 2118 1025 2121
rect 1677 2118 1678 2122
rect 1746 2118 1747 2122
rect 1941 2118 1942 2122
rect 3146 2118 3148 2122
rect 992 2103 994 2107
rect 998 2103 1001 2107
rect 1005 2103 1008 2107
rect 2024 2103 2026 2107
rect 2030 2103 2033 2107
rect 2037 2103 2040 2107
rect 3040 2103 3042 2107
rect 3046 2103 3049 2107
rect 3053 2103 3056 2107
rect 1789 2088 1790 2092
rect 1962 2088 1963 2092
rect 2013 2088 2014 2092
rect 3170 2088 3172 2092
rect 3213 2088 3214 2092
rect 14 2058 33 2061
rect 62 2061 65 2071
rect 222 2068 233 2071
rect 718 2068 729 2071
rect 798 2068 809 2071
rect 846 2068 857 2071
rect 1254 2068 1262 2071
rect 1350 2068 1361 2071
rect 1710 2068 1718 2071
rect 1798 2068 1817 2071
rect 2046 2071 2049 2081
rect 2554 2078 2569 2081
rect 2734 2072 2737 2081
rect 2026 2068 2049 2071
rect 2054 2068 2062 2071
rect 2490 2068 2497 2071
rect 2538 2068 2577 2071
rect 2686 2068 2705 2071
rect 2822 2071 2825 2081
rect 3250 2078 3257 2081
rect 2806 2068 2825 2071
rect 2838 2068 2865 2071
rect 2930 2068 2945 2071
rect 2998 2068 3009 2071
rect 3058 2068 3065 2071
rect 3082 2068 3089 2071
rect 3342 2068 3353 2071
rect 718 2062 721 2068
rect 3350 2062 3353 2068
rect 50 2058 65 2061
rect 202 2058 209 2061
rect 410 2058 425 2061
rect 470 2058 489 2061
rect 582 2058 590 2061
rect 634 2058 646 2061
rect 678 2058 697 2061
rect 810 2058 817 2061
rect 878 2058 897 2061
rect 954 2058 969 2061
rect 978 2058 1017 2061
rect 1062 2058 1081 2061
rect 1126 2058 1134 2061
rect 1158 2058 1174 2061
rect 1226 2058 1241 2061
rect 1294 2058 1313 2061
rect 1450 2058 1462 2061
rect 1506 2058 1529 2061
rect 1558 2058 1566 2061
rect 1670 2058 1689 2061
rect 1766 2058 1774 2061
rect 2470 2058 2489 2061
rect 2662 2058 2670 2061
rect 2990 2058 2998 2061
rect 3050 2058 3057 2061
rect 3246 2058 3257 2061
rect 3362 2058 3369 2061
rect 3374 2058 3393 2061
rect 30 2048 33 2058
rect 422 2048 425 2058
rect 470 2048 473 2058
rect 694 2048 697 2058
rect 878 2048 881 2058
rect 1062 2048 1065 2058
rect 1134 2048 1153 2051
rect 1158 2048 1161 2058
rect 1310 2048 1313 2058
rect 1478 2048 1497 2051
rect 1582 2048 1601 2051
rect 1686 2048 1689 2058
rect 1746 2048 1753 2051
rect 1882 2048 1889 2051
rect 2694 2048 2702 2051
rect 2986 2048 2990 2052
rect 1862 2042 1866 2044
rect 1018 2038 1019 2042
rect 2364 2038 2366 2042
rect 2762 2038 2769 2041
rect 3180 2038 3182 2042
rect 3290 2038 3292 2042
rect 3542 2038 3558 2041
rect 45 2018 46 2022
rect 98 2018 99 2022
rect 178 2018 179 2022
rect 261 2018 262 2022
rect 322 2018 323 2022
rect 530 2018 531 2022
rect 738 2018 739 2022
rect 770 2018 771 2022
rect 818 2018 819 2022
rect 866 2018 867 2022
rect 941 2018 942 2022
rect 1050 2018 1051 2022
rect 1178 2018 1179 2022
rect 1213 2018 1214 2022
rect 1370 2018 1371 2022
rect 1466 2018 1467 2022
rect 1546 2018 1547 2022
rect 1613 2018 1614 2022
rect 1730 2018 1731 2022
rect 1845 2018 1846 2022
rect 2197 2018 2198 2022
rect 3242 2018 3243 2022
rect 3509 2018 3510 2022
rect 480 2003 482 2007
rect 486 2003 489 2007
rect 493 2003 496 2007
rect 1512 2003 1514 2007
rect 1518 2003 1521 2007
rect 1525 2003 1528 2007
rect 2536 2003 2538 2007
rect 2542 2003 2545 2007
rect 2549 2003 2552 2007
rect 658 1988 659 1992
rect 1373 1988 1374 1992
rect 1405 1988 1406 1992
rect 1602 1988 1603 1992
rect 2042 1988 2043 1992
rect 2170 1988 2171 1992
rect 2386 1988 2387 1992
rect 2570 1988 2571 1992
rect 2994 1988 2995 1992
rect 1726 1972 1729 1981
rect 74 1968 82 1971
rect 770 1968 771 1972
rect 894 1968 914 1971
rect 1021 1968 1022 1972
rect 1106 1968 1107 1972
rect 2202 1968 2209 1971
rect 3430 1968 3441 1971
rect 3430 1962 3433 1968
rect 30 1958 49 1961
rect 54 1958 65 1961
rect 110 1951 113 1961
rect 438 1958 457 1961
rect 974 1958 1009 1961
rect 98 1948 113 1951
rect 138 1948 145 1951
rect 262 1948 270 1951
rect 314 1948 321 1951
rect 354 1948 361 1951
rect 470 1948 478 1951
rect 518 1948 526 1951
rect 674 1948 681 1951
rect 838 1948 846 1951
rect 850 1948 865 1951
rect 1118 1951 1121 1961
rect 1174 1951 1177 1961
rect 1082 1948 1105 1951
rect 1118 1948 1137 1951
rect 1158 1948 1177 1951
rect 1230 1951 1233 1961
rect 1614 1958 1625 1961
rect 2146 1958 2153 1961
rect 2186 1958 2193 1961
rect 3250 1958 3254 1962
rect 3438 1958 3449 1961
rect 1210 1948 1217 1951
rect 1230 1948 1249 1951
rect 1330 1948 1337 1951
rect 1554 1948 1561 1951
rect 1582 1948 1598 1951
rect 2006 1948 2038 1951
rect 2534 1948 2550 1951
rect 2846 1951 2849 1958
rect 3422 1956 3426 1958
rect 2838 1948 2849 1951
rect 3190 1948 3209 1951
rect 3242 1948 3249 1951
rect 262 1938 265 1948
rect 358 1938 361 1948
rect 558 1938 566 1941
rect 642 1938 649 1941
rect 698 1938 705 1941
rect 1146 1938 1153 1941
rect 1258 1938 1265 1941
rect 1442 1938 1457 1941
rect 1658 1938 1665 1941
rect 1806 1938 1814 1941
rect 2638 1941 2641 1948
rect 3478 1942 3481 1951
rect 2630 1938 2641 1941
rect 3022 1938 3038 1941
rect 3274 1938 3281 1941
rect 3314 1938 3321 1941
rect 3542 1938 3558 1941
rect 157 1928 158 1932
rect 206 1928 217 1931
rect 1982 1928 2001 1931
rect 2086 1931 2089 1938
rect 2070 1928 2089 1931
rect 2894 1928 2905 1931
rect 3422 1931 3426 1933
rect 3422 1928 3433 1931
rect 370 1918 371 1922
rect 389 1918 390 1922
rect 741 1918 742 1922
rect 954 1918 955 1922
rect 1045 1918 1046 1922
rect 992 1903 994 1907
rect 998 1903 1001 1907
rect 1005 1903 1008 1907
rect 2024 1903 2026 1907
rect 2030 1903 2033 1907
rect 2037 1903 2040 1907
rect 3040 1903 3042 1907
rect 3046 1903 3049 1907
rect 3053 1903 3056 1907
rect 1330 1888 1331 1892
rect 1661 1888 1662 1892
rect 1786 1888 1787 1892
rect 1146 1878 1147 1882
rect 2042 1878 2057 1881
rect 2534 1878 2564 1881
rect 2766 1878 2782 1881
rect 3026 1878 3038 1881
rect 10 1868 17 1871
rect 126 1868 137 1871
rect 198 1868 209 1871
rect 334 1868 342 1871
rect 406 1868 422 1871
rect 734 1868 742 1871
rect 894 1868 913 1871
rect 1018 1868 1025 1871
rect 1218 1868 1233 1871
rect 1382 1868 1409 1871
rect 1522 1868 1537 1871
rect 1542 1868 1561 1871
rect 1742 1868 1750 1871
rect 1782 1868 1801 1871
rect 1902 1868 1929 1871
rect 1974 1868 1982 1871
rect 2022 1868 2046 1871
rect 2070 1868 2086 1871
rect 2342 1868 2350 1871
rect 2362 1868 2369 1871
rect 2622 1868 2633 1871
rect 2670 1868 2678 1871
rect 2806 1868 2825 1871
rect 2866 1868 2873 1871
rect 2910 1868 2918 1871
rect 2994 1868 3001 1871
rect 3046 1868 3073 1871
rect 158 1858 177 1861
rect 258 1858 281 1861
rect 286 1858 294 1861
rect 298 1858 305 1861
rect 406 1858 430 1861
rect 538 1858 545 1861
rect 622 1858 641 1861
rect 702 1858 721 1861
rect 786 1858 793 1861
rect 854 1858 862 1861
rect 1226 1858 1233 1861
rect 1266 1858 1273 1861
rect 1682 1858 1689 1861
rect 1694 1858 1702 1861
rect 1802 1858 1809 1861
rect 1814 1858 1822 1861
rect 1854 1858 1862 1861
rect 2118 1858 2121 1868
rect 2622 1862 2625 1868
rect 2382 1858 2402 1861
rect 2662 1861 2665 1868
rect 3070 1862 3073 1868
rect 2654 1858 2665 1861
rect 2714 1858 2721 1861
rect 3102 1858 3110 1861
rect 3134 1858 3142 1861
rect 3346 1858 3353 1861
rect 3406 1858 3414 1861
rect 3530 1858 3537 1861
rect 174 1848 177 1858
rect 638 1848 641 1858
rect 718 1852 721 1858
rect 746 1848 753 1851
rect 862 1848 881 1851
rect 886 1848 897 1851
rect 934 1848 953 1851
rect 1054 1848 1073 1851
rect 1078 1848 1097 1851
rect 3204 1848 3206 1852
rect 1070 1842 1074 1844
rect 726 1838 734 1841
rect 1290 1838 1291 1842
rect 2962 1838 2964 1842
rect 3550 1838 3558 1841
rect 61 1818 62 1822
rect 581 1818 582 1822
rect 653 1818 654 1822
rect 701 1818 702 1822
rect 1194 1818 1195 1822
rect 1450 1818 1451 1822
rect 2722 1818 2723 1822
rect 480 1803 482 1807
rect 486 1803 489 1807
rect 493 1803 496 1807
rect 1512 1803 1514 1807
rect 1518 1803 1521 1807
rect 1525 1803 1528 1807
rect 2536 1803 2538 1807
rect 2542 1803 2545 1807
rect 2549 1803 2552 1807
rect 1197 1788 1198 1792
rect 1490 1788 1491 1792
rect 1602 1788 1603 1792
rect 1786 1788 1787 1792
rect 2258 1788 2259 1792
rect 2677 1788 2678 1792
rect 3154 1788 3155 1792
rect 3282 1788 3283 1792
rect 3397 1788 3398 1792
rect 722 1778 723 1782
rect 1133 1778 1134 1782
rect 1725 1778 1726 1782
rect 1826 1778 1827 1782
rect 1925 1778 1926 1782
rect 2722 1768 2729 1771
rect 82 1748 94 1751
rect 598 1748 606 1751
rect 650 1748 657 1751
rect 678 1751 681 1761
rect 826 1758 833 1761
rect 838 1758 857 1761
rect 678 1748 697 1751
rect 714 1748 721 1751
rect 770 1748 785 1751
rect 870 1748 878 1751
rect 882 1748 897 1751
rect 1062 1751 1065 1761
rect 1102 1758 1121 1761
rect 1286 1761 1289 1768
rect 1286 1758 1297 1761
rect 1502 1758 1518 1761
rect 1538 1758 1542 1762
rect 3025 1758 3033 1762
rect 1046 1748 1065 1751
rect 1134 1748 1150 1751
rect 1270 1748 1278 1751
rect 1318 1748 1345 1751
rect 1514 1748 1537 1751
rect 1682 1748 1689 1751
rect 1746 1748 1753 1751
rect 1758 1748 1785 1751
rect 1874 1748 1881 1751
rect 2130 1748 2150 1751
rect 2718 1751 2721 1758
rect 3030 1752 3033 1758
rect 2710 1748 2721 1751
rect 2758 1748 2769 1751
rect 2870 1748 2878 1751
rect 3166 1751 3169 1758
rect 3166 1748 3177 1751
rect 3266 1748 3281 1751
rect 3334 1748 3350 1751
rect 78 1738 81 1748
rect 198 1741 201 1748
rect 198 1738 209 1741
rect 326 1738 345 1741
rect 478 1738 494 1741
rect 550 1738 577 1741
rect 654 1738 657 1748
rect 766 1741 769 1748
rect 758 1738 769 1741
rect 986 1738 1009 1741
rect 1582 1738 1585 1748
rect 1734 1738 1742 1741
rect 1806 1738 1814 1741
rect 1870 1738 1881 1741
rect 1934 1738 1953 1741
rect 1962 1738 1969 1741
rect 2142 1738 2150 1741
rect 2202 1738 2209 1741
rect 2238 1738 2249 1741
rect 2518 1738 2553 1741
rect 2846 1738 2865 1741
rect 2886 1738 2913 1741
rect 2926 1738 2974 1741
rect 3046 1738 3062 1741
rect 3118 1738 3137 1741
rect 38 1732 41 1738
rect 958 1732 961 1738
rect 1878 1732 1881 1738
rect 3206 1732 3209 1738
rect 3470 1732 3474 1734
rect 38 1728 46 1732
rect 954 1728 961 1732
rect 1234 1728 1235 1732
rect 2190 1728 2201 1731
rect 2702 1728 2721 1731
rect 3206 1728 3214 1732
rect 3242 1728 3249 1731
rect 3558 1728 3561 1738
rect 130 1718 131 1722
rect 522 1718 523 1722
rect 618 1718 619 1722
rect 2014 1718 2030 1721
rect 992 1703 994 1707
rect 998 1703 1001 1707
rect 1005 1703 1008 1707
rect 2024 1703 2026 1707
rect 2030 1703 2033 1707
rect 2037 1703 2040 1707
rect 3040 1703 3042 1707
rect 3046 1703 3049 1707
rect 3053 1703 3056 1707
rect 29 1688 30 1692
rect 1461 1688 1462 1692
rect 1502 1688 1518 1691
rect 2322 1688 2323 1692
rect 2613 1688 2614 1692
rect 2669 1688 2670 1692
rect 78 1668 86 1671
rect 126 1668 145 1671
rect 614 1671 617 1681
rect 646 1678 654 1681
rect 1094 1678 1110 1681
rect 1786 1678 1787 1682
rect 1934 1672 1937 1681
rect 2146 1678 2153 1681
rect 2970 1678 2977 1681
rect 3342 1678 3353 1681
rect 590 1668 601 1671
rect 614 1668 622 1671
rect 638 1668 646 1671
rect 1646 1668 1657 1671
rect 1666 1668 1673 1671
rect 1750 1668 1758 1671
rect 1910 1668 1918 1671
rect 1938 1668 1945 1671
rect 1970 1668 1977 1671
rect 2006 1668 2025 1671
rect 2070 1668 2078 1671
rect 2582 1671 2585 1678
rect 3342 1672 3345 1678
rect 3358 1672 3361 1681
rect 2582 1668 2593 1671
rect 2754 1668 2761 1671
rect 2782 1668 2793 1671
rect 2934 1668 2942 1671
rect 3370 1668 3377 1671
rect 3526 1668 3545 1671
rect 598 1662 601 1668
rect 2782 1662 2785 1668
rect 10 1658 17 1661
rect 174 1658 193 1661
rect 286 1658 294 1661
rect 318 1658 334 1661
rect 462 1658 494 1661
rect 542 1658 558 1661
rect 774 1658 793 1661
rect 814 1658 833 1661
rect 850 1658 865 1661
rect 906 1658 913 1661
rect 950 1658 966 1661
rect 1046 1658 1054 1661
rect 1070 1658 1078 1661
rect 1138 1658 1153 1661
rect 1178 1658 1185 1661
rect 2030 1658 2038 1661
rect 2390 1658 2417 1661
rect 2518 1658 2526 1661
rect 2842 1658 2849 1661
rect 2938 1658 2945 1661
rect 3022 1658 3033 1661
rect 3126 1658 3134 1661
rect 3154 1658 3161 1661
rect 3206 1658 3214 1661
rect 3286 1658 3294 1661
rect 3334 1658 3342 1661
rect 3406 1658 3414 1661
rect 3454 1661 3457 1668
rect 3454 1658 3465 1661
rect 190 1648 193 1658
rect 506 1648 510 1652
rect 542 1648 545 1658
rect 774 1648 777 1658
rect 830 1648 833 1658
rect 862 1648 865 1658
rect 938 1648 945 1651
rect 950 1648 953 1658
rect 1298 1648 1305 1651
rect 1314 1648 1318 1652
rect 1502 1648 1518 1651
rect 1634 1648 1638 1652
rect 2526 1648 2542 1651
rect 3030 1648 3046 1651
rect 3318 1648 3326 1651
rect 3402 1648 3406 1652
rect 90 1638 97 1641
rect 205 1638 206 1642
rect 530 1638 537 1641
rect 733 1638 734 1642
rect 870 1638 878 1641
rect 357 1628 358 1632
rect 69 1618 70 1622
rect 285 1618 286 1622
rect 698 1618 699 1622
rect 762 1618 763 1622
rect 1029 1618 1030 1622
rect 1069 1618 1070 1622
rect 1154 1618 1155 1622
rect 1925 1618 1926 1622
rect 2485 1618 2486 1622
rect 2730 1618 2731 1622
rect 3074 1618 3075 1622
rect 480 1603 482 1607
rect 486 1603 489 1607
rect 493 1603 496 1607
rect 1512 1603 1514 1607
rect 1518 1603 1521 1607
rect 1525 1603 1528 1607
rect 2536 1603 2538 1607
rect 2542 1603 2545 1607
rect 2549 1603 2552 1607
rect 1242 1588 1243 1592
rect 1434 1588 1435 1592
rect 1597 1588 1598 1592
rect 1957 1588 1958 1592
rect 2069 1588 2070 1592
rect 2213 1588 2214 1592
rect 2853 1588 2854 1592
rect 3373 1588 3374 1592
rect 306 1568 307 1572
rect 413 1568 414 1572
rect 925 1568 926 1572
rect 2013 1568 2014 1572
rect 2542 1568 2550 1571
rect 2746 1568 2761 1571
rect 3550 1568 3558 1571
rect 134 1548 142 1551
rect 242 1548 249 1551
rect 322 1548 329 1551
rect 418 1548 433 1551
rect 518 1551 521 1561
rect 518 1548 537 1551
rect 546 1548 553 1551
rect 558 1548 566 1551
rect 574 1548 582 1551
rect 638 1551 641 1561
rect 626 1548 641 1551
rect 666 1548 673 1551
rect 782 1551 785 1561
rect 986 1558 993 1561
rect 1062 1552 1065 1561
rect 766 1548 785 1551
rect 902 1548 910 1551
rect 998 1548 1022 1551
rect 1082 1548 1089 1551
rect 1142 1551 1145 1561
rect 1198 1558 1217 1561
rect 1126 1548 1145 1551
rect 1178 1548 1185 1551
rect 1234 1548 1241 1551
rect 1318 1551 1321 1568
rect 1302 1548 1321 1551
rect 1334 1552 1337 1561
rect 1362 1548 1377 1551
rect 1382 1548 1398 1551
rect 1418 1548 1433 1551
rect 1482 1548 1489 1551
rect 1738 1548 1745 1551
rect 1818 1548 1833 1551
rect 2034 1548 2057 1551
rect 2198 1551 2201 1561
rect 2182 1548 2201 1551
rect 2278 1548 2286 1551
rect 58 1538 65 1541
rect 110 1538 118 1541
rect 430 1538 433 1548
rect 662 1538 665 1548
rect 694 1541 697 1548
rect 750 1541 753 1548
rect 678 1538 697 1541
rect 742 1538 753 1541
rect 834 1538 849 1541
rect 1094 1541 1097 1548
rect 1094 1538 1105 1541
rect 1478 1538 1489 1541
rect 1494 1538 1518 1541
rect 1642 1538 1649 1541
rect 1790 1538 1809 1541
rect 2322 1538 2329 1541
rect 2414 1541 2417 1548
rect 2710 1542 2713 1551
rect 3034 1548 3057 1551
rect 3082 1548 3089 1551
rect 3290 1548 3297 1551
rect 2414 1538 2425 1541
rect 2562 1538 2577 1541
rect 2682 1538 2697 1541
rect 2914 1538 2926 1541
rect 2942 1538 2950 1541
rect 3234 1538 3242 1541
rect 3358 1538 3366 1541
rect 3418 1538 3425 1541
rect 154 1528 158 1532
rect 1262 1531 1265 1538
rect 1486 1532 1489 1538
rect 1262 1528 1273 1531
rect 1686 1528 1694 1531
rect 1770 1528 1777 1531
rect 1918 1531 1921 1538
rect 1918 1528 1929 1531
rect 1934 1528 1945 1531
rect 2342 1528 2353 1531
rect 2710 1528 2729 1531
rect 3382 1528 3393 1531
rect 50 1518 51 1522
rect 74 1518 75 1522
rect 186 1518 187 1522
rect 442 1518 443 1522
rect 826 1518 827 1522
rect 978 1518 979 1522
rect 1522 1518 1529 1521
rect 992 1503 994 1507
rect 998 1503 1001 1507
rect 1005 1503 1008 1507
rect 2024 1503 2026 1507
rect 2030 1503 2033 1507
rect 2037 1503 2040 1507
rect 3040 1503 3042 1507
rect 3046 1503 3049 1507
rect 3053 1503 3056 1507
rect 674 1488 675 1492
rect 1133 1488 1134 1492
rect 1477 1488 1478 1492
rect 1538 1488 1545 1491
rect 1890 1488 1891 1492
rect 2077 1488 2078 1492
rect 2538 1488 2553 1491
rect 338 1478 345 1481
rect 1518 1478 1534 1481
rect 14 1468 25 1471
rect 462 1462 465 1471
rect 714 1468 721 1471
rect 766 1462 769 1471
rect 806 1468 817 1471
rect 854 1468 865 1471
rect 1282 1468 1297 1471
rect 1406 1468 1414 1471
rect 1454 1468 1470 1471
rect 1582 1471 1585 1481
rect 1638 1478 1646 1481
rect 2510 1478 2521 1481
rect 3022 1472 3025 1481
rect 3454 1478 3465 1481
rect 3542 1478 3550 1482
rect 3454 1472 3457 1478
rect 3542 1472 3545 1478
rect 1562 1468 1569 1471
rect 1582 1468 1590 1471
rect 1698 1468 1713 1471
rect 26 1458 33 1461
rect 38 1458 65 1461
rect 106 1458 113 1461
rect 134 1458 153 1461
rect 406 1458 433 1461
rect 514 1458 521 1461
rect 630 1458 649 1461
rect 734 1458 750 1461
rect 886 1458 905 1461
rect 958 1458 974 1461
rect 1046 1458 1062 1461
rect 1114 1458 1121 1461
rect 1326 1458 1342 1461
rect 1490 1458 1505 1461
rect 1766 1461 1769 1468
rect 1758 1458 1769 1461
rect 1810 1458 1817 1461
rect 1822 1458 1849 1461
rect 2062 1458 2070 1461
rect 2142 1458 2150 1461
rect 2230 1458 2238 1461
rect 2270 1458 2278 1461
rect 2302 1458 2310 1461
rect 2382 1458 2393 1461
rect 2446 1458 2454 1461
rect 2478 1461 2481 1471
rect 2562 1468 2577 1471
rect 2646 1468 2665 1471
rect 2694 1468 2705 1471
rect 2790 1468 2809 1471
rect 2986 1468 3001 1471
rect 3074 1468 3082 1471
rect 3198 1468 3209 1471
rect 3482 1468 3489 1471
rect 2662 1462 2665 1468
rect 2478 1458 2486 1461
rect 2490 1458 2497 1461
rect 2522 1458 2529 1461
rect 2562 1458 2569 1461
rect 2726 1458 2737 1461
rect 2758 1458 2766 1461
rect 2814 1458 2838 1461
rect 2894 1458 2902 1461
rect 2982 1458 2990 1461
rect 3178 1458 3185 1461
rect 3222 1458 3230 1461
rect 3262 1458 3270 1461
rect 3534 1458 3553 1461
rect 86 1448 94 1451
rect 150 1448 153 1458
rect 630 1448 633 1458
rect 734 1448 737 1458
rect 886 1448 889 1458
rect 2726 1452 2729 1458
rect 966 1448 985 1451
rect 990 1448 1006 1451
rect 2670 1448 2678 1451
rect 3218 1448 3222 1452
rect 3330 1448 3337 1451
rect 237 1438 238 1442
rect 618 1438 619 1442
rect 874 1438 875 1442
rect 922 1438 929 1441
rect 1794 1438 1801 1441
rect 3014 1438 3022 1441
rect 66 1428 67 1432
rect 1085 1428 1086 1432
rect 1173 1428 1174 1432
rect 34 1418 35 1422
rect 165 1418 166 1422
rect 197 1418 198 1422
rect 277 1418 278 1422
rect 373 1418 374 1422
rect 533 1418 534 1422
rect 581 1418 582 1422
rect 1914 1418 1915 1422
rect 1949 1418 1950 1422
rect 1973 1418 1974 1422
rect 2378 1418 2379 1422
rect 2781 1418 2782 1422
rect 480 1403 482 1407
rect 486 1403 489 1407
rect 493 1403 496 1407
rect 1512 1403 1514 1407
rect 1518 1403 1521 1407
rect 1525 1403 1528 1407
rect 2536 1403 2538 1407
rect 2542 1403 2545 1407
rect 2549 1403 2552 1407
rect 509 1388 510 1392
rect 1282 1388 1283 1392
rect 1314 1388 1315 1392
rect 1450 1388 1451 1392
rect 2274 1388 2275 1392
rect 2866 1388 2867 1392
rect 3148 1388 3150 1392
rect 3402 1388 3404 1392
rect 3453 1388 3454 1392
rect 2989 1378 2990 1382
rect 610 1368 611 1372
rect 1738 1368 1753 1371
rect 2286 1368 2297 1371
rect 2514 1368 2521 1371
rect 158 1358 166 1361
rect 206 1358 214 1361
rect 430 1358 441 1361
rect 490 1358 497 1361
rect 622 1358 641 1361
rect 1226 1358 1230 1362
rect 1482 1358 1486 1362
rect 1562 1358 1569 1361
rect 1882 1358 1889 1361
rect 1894 1358 1902 1361
rect 438 1352 441 1358
rect 78 1348 86 1351
rect 510 1348 526 1351
rect 738 1348 753 1351
rect 822 1348 830 1351
rect 1206 1348 1214 1351
rect 1254 1348 1281 1351
rect 1298 1348 1305 1351
rect 1422 1348 1449 1351
rect 1526 1351 1529 1358
rect 1510 1348 1529 1351
rect 1550 1348 1566 1351
rect 1594 1348 1601 1351
rect 1606 1348 1633 1351
rect 1802 1348 1809 1351
rect 1850 1348 1865 1351
rect 78 1338 81 1348
rect 126 1338 134 1341
rect 278 1338 289 1341
rect 366 1338 374 1341
rect 594 1338 601 1341
rect 650 1338 657 1341
rect 674 1338 681 1341
rect 762 1338 769 1341
rect 846 1338 857 1341
rect 1086 1338 1102 1341
rect 1142 1338 1161 1341
rect 1302 1338 1305 1348
rect 1350 1341 1353 1348
rect 2062 1342 2065 1351
rect 2398 1348 2417 1351
rect 1342 1338 1353 1341
rect 1522 1338 1542 1341
rect 1706 1338 1713 1341
rect 1794 1338 1801 1341
rect 1846 1338 1854 1341
rect 1946 1338 1953 1341
rect 2234 1338 2241 1341
rect 2470 1341 2473 1351
rect 2586 1348 2593 1351
rect 2658 1348 2665 1351
rect 3198 1351 3201 1361
rect 3150 1348 3185 1351
rect 3198 1348 3217 1351
rect 2438 1338 2457 1341
rect 2470 1338 2489 1341
rect 3006 1341 3009 1348
rect 3006 1338 3017 1341
rect 3246 1338 3265 1341
rect 3534 1341 3537 1348
rect 3526 1338 3537 1341
rect 1158 1328 1161 1338
rect 2006 1328 2014 1331
rect 2018 1328 2033 1331
rect 2110 1328 2121 1331
rect 2310 1328 2329 1331
rect 2454 1328 2457 1338
rect 2462 1328 2470 1331
rect 2782 1328 2793 1331
rect 3262 1328 3265 1338
rect 2110 1322 2113 1328
rect 13 1318 14 1322
rect 37 1318 38 1322
rect 98 1318 99 1322
rect 154 1318 155 1322
rect 178 1318 179 1322
rect 386 1318 387 1322
rect 470 1318 486 1321
rect 581 1318 582 1322
rect 778 1318 779 1322
rect 970 1318 971 1322
rect 1037 1318 1038 1322
rect 2538 1318 2553 1321
rect 992 1303 994 1307
rect 998 1303 1001 1307
rect 1005 1303 1008 1307
rect 2024 1303 2026 1307
rect 2030 1303 2033 1307
rect 2037 1303 2040 1307
rect 3040 1303 3042 1307
rect 3046 1303 3049 1307
rect 3053 1303 3056 1307
rect 61 1288 62 1292
rect 1893 1288 1894 1292
rect 2197 1288 2198 1292
rect 2542 1288 2558 1291
rect 2794 1288 2795 1292
rect 2845 1288 2846 1292
rect 3084 1288 3086 1292
rect 746 1278 753 1281
rect 1002 1278 1014 1281
rect 1026 1278 1033 1281
rect 110 1268 121 1271
rect 150 1268 158 1271
rect 202 1268 209 1271
rect 278 1268 286 1271
rect 306 1268 313 1271
rect 390 1268 401 1271
rect 530 1268 537 1271
rect 618 1268 625 1271
rect 834 1268 841 1271
rect 990 1268 1022 1271
rect 398 1262 401 1268
rect 102 1258 110 1261
rect 174 1258 182 1261
rect 458 1258 473 1261
rect 574 1258 593 1261
rect 590 1252 593 1258
rect 610 1258 617 1261
rect 818 1258 833 1261
rect 918 1258 942 1261
rect 1010 1258 1025 1261
rect 1118 1261 1121 1281
rect 1578 1278 1585 1281
rect 1758 1278 1766 1281
rect 1842 1278 1849 1282
rect 2042 1278 2049 1281
rect 1846 1272 1849 1278
rect 1154 1268 1161 1271
rect 1178 1268 1193 1271
rect 1394 1268 1401 1271
rect 1486 1268 1510 1271
rect 1118 1258 1126 1261
rect 1354 1261 1361 1264
rect 1470 1258 1481 1261
rect 1534 1258 1542 1261
rect 1606 1258 1625 1261
rect 1654 1261 1657 1271
rect 1902 1262 1905 1271
rect 1942 1268 1961 1271
rect 1990 1268 2006 1271
rect 2062 1268 2081 1271
rect 2182 1268 2201 1271
rect 2286 1268 2294 1271
rect 2342 1268 2361 1271
rect 2546 1268 2577 1271
rect 2698 1268 2705 1271
rect 2766 1268 2793 1271
rect 2806 1268 2825 1271
rect 3006 1268 3014 1271
rect 3106 1268 3113 1271
rect 3302 1271 3305 1281
rect 3298 1268 3305 1271
rect 3390 1268 3398 1271
rect 1650 1258 1657 1261
rect 1838 1258 1857 1261
rect 2142 1258 2158 1261
rect 2174 1258 2190 1261
rect 2210 1258 2225 1261
rect 2278 1258 2289 1261
rect 2554 1258 2569 1261
rect 2586 1258 2601 1261
rect 2878 1258 2886 1261
rect 2898 1258 2905 1261
rect 2942 1258 2961 1261
rect 3114 1258 3121 1261
rect 3126 1258 3137 1261
rect 3142 1258 3166 1261
rect 3174 1258 3190 1261
rect 3230 1258 3238 1261
rect 3390 1258 3409 1261
rect 186 1248 193 1251
rect 606 1248 609 1258
rect 758 1248 769 1251
rect 914 1248 918 1252
rect 1506 1248 1521 1251
rect 1530 1248 1534 1252
rect 1622 1248 1625 1258
rect 1782 1248 1801 1251
rect 1854 1248 1857 1258
rect 2286 1252 2289 1258
rect 2942 1252 2945 1258
rect 3126 1252 3129 1258
rect 1929 1248 1934 1252
rect 2266 1248 2273 1251
rect 2874 1248 2878 1252
rect 2990 1248 3001 1251
rect 3186 1248 3193 1251
rect 3210 1248 3217 1251
rect 3282 1248 3289 1251
rect 3390 1248 3393 1258
rect 238 1238 246 1241
rect 421 1238 422 1242
rect 1245 1238 1246 1242
rect 1558 1238 1566 1241
rect 1813 1228 1814 1232
rect 101 1218 102 1222
rect 322 1218 323 1222
rect 685 1218 686 1222
rect 781 1218 782 1222
rect 957 1218 958 1222
rect 1637 1218 1638 1222
rect 2038 1221 2041 1228
rect 2038 1218 2049 1221
rect 2173 1218 2174 1222
rect 480 1203 482 1207
rect 486 1203 489 1207
rect 493 1203 496 1207
rect 1512 1203 1514 1207
rect 1518 1203 1521 1207
rect 1525 1203 1528 1207
rect 2536 1203 2538 1207
rect 2542 1203 2545 1207
rect 2549 1203 2552 1207
rect 18 1188 19 1192
rect 146 1188 147 1192
rect 237 1188 238 1192
rect 565 1188 566 1192
rect 1026 1188 1027 1192
rect 1077 1188 1078 1192
rect 1277 1188 1278 1192
rect 1314 1188 1315 1192
rect 1437 1188 1438 1192
rect 1562 1188 1563 1192
rect 1642 1188 1643 1192
rect 1861 1188 1862 1192
rect 2542 1188 2558 1191
rect 2917 1188 2918 1192
rect 2941 1188 2942 1192
rect 2970 1188 2971 1192
rect 3018 1188 3019 1192
rect 3054 1188 3070 1191
rect 402 1178 403 1182
rect 1354 1178 1355 1182
rect 2869 1178 2870 1182
rect 293 1168 294 1172
rect 1198 1168 1209 1171
rect 1469 1168 1470 1172
rect 3410 1168 3425 1171
rect 3558 1171 3561 1178
rect 3550 1168 3561 1171
rect 1206 1162 1209 1168
rect 186 1158 193 1161
rect 438 1158 446 1161
rect 34 1148 49 1151
rect 194 1148 201 1151
rect 450 1148 457 1151
rect 474 1148 497 1151
rect 526 1148 534 1151
rect 670 1148 686 1151
rect 702 1151 705 1161
rect 702 1148 718 1151
rect 782 1151 785 1161
rect 782 1148 801 1151
rect 850 1148 857 1151
rect 246 1138 265 1141
rect 382 1138 390 1141
rect 598 1138 606 1141
rect 694 1138 702 1141
rect 878 1141 881 1148
rect 870 1138 881 1141
rect 894 1141 897 1151
rect 1042 1148 1049 1151
rect 1090 1148 1105 1151
rect 1210 1148 1217 1151
rect 1222 1148 1238 1151
rect 1262 1151 1265 1161
rect 1366 1158 1385 1161
rect 1686 1152 1689 1161
rect 2030 1158 2038 1161
rect 1246 1148 1265 1151
rect 1326 1148 1342 1151
rect 1522 1148 1550 1151
rect 1658 1148 1673 1151
rect 1886 1151 1890 1152
rect 1874 1148 1890 1151
rect 1914 1148 1921 1151
rect 1926 1148 1934 1151
rect 2238 1148 2249 1151
rect 2282 1148 2297 1151
rect 2470 1148 2481 1151
rect 2750 1148 2766 1151
rect 2854 1151 2857 1161
rect 2838 1148 2857 1151
rect 2870 1148 2889 1151
rect 2922 1148 2937 1151
rect 2954 1148 2969 1151
rect 3054 1148 3078 1151
rect 3106 1148 3113 1151
rect 3142 1151 3145 1161
rect 3142 1148 3158 1151
rect 3190 1148 3198 1151
rect 3234 1148 3246 1151
rect 2246 1142 2249 1148
rect 894 1138 913 1141
rect 966 1138 974 1141
rect 1086 1138 1094 1141
rect 1234 1138 1241 1141
rect 1518 1138 1526 1141
rect 1614 1138 1622 1141
rect 1738 1138 1745 1141
rect 1938 1138 1945 1141
rect 2150 1138 2158 1141
rect 2282 1138 2289 1141
rect 2310 1138 2329 1141
rect 2398 1138 2406 1141
rect 2598 1138 2606 1141
rect 2630 1138 2638 1141
rect 2694 1138 2702 1141
rect 2758 1138 2777 1141
rect 2950 1138 2958 1141
rect 2994 1138 3001 1141
rect 3086 1138 3102 1141
rect 3134 1138 3142 1141
rect 3198 1138 3217 1141
rect 3226 1138 3241 1141
rect 3262 1138 3273 1141
rect 3342 1138 3350 1141
rect 350 1128 361 1131
rect 925 1128 926 1132
rect 1054 1128 1057 1138
rect 2562 1128 2569 1131
rect 2950 1128 2953 1138
rect 3182 1131 3185 1138
rect 3098 1128 3105 1131
rect 3174 1128 3185 1131
rect 3198 1128 3201 1138
rect 122 1118 123 1122
rect 434 1118 435 1122
rect 546 1118 547 1122
rect 589 1118 590 1122
rect 733 1118 734 1122
rect 962 1118 963 1122
rect 986 1118 987 1122
rect 1117 1118 1118 1122
rect 1818 1118 1819 1122
rect 2490 1118 2491 1122
rect 3300 1118 3302 1122
rect 992 1103 994 1107
rect 998 1103 1001 1107
rect 1005 1103 1008 1107
rect 2024 1103 2026 1107
rect 2030 1103 2033 1107
rect 2037 1103 2040 1107
rect 3040 1103 3042 1107
rect 3046 1103 3049 1107
rect 3053 1103 3056 1107
rect 1157 1088 1158 1092
rect 3213 1088 3214 1092
rect 3237 1088 3238 1092
rect 1074 1078 1081 1081
rect 1406 1078 1417 1081
rect 1466 1078 1473 1081
rect 1878 1078 1889 1081
rect 2014 1078 2049 1081
rect 1886 1072 1889 1078
rect 30 1068 41 1071
rect 58 1068 65 1071
rect 94 1068 105 1071
rect 222 1068 238 1071
rect 158 1058 166 1061
rect 190 1058 198 1061
rect 246 1058 265 1061
rect 294 1061 297 1071
rect 290 1058 297 1061
rect 310 1058 329 1061
rect 358 1058 374 1061
rect 470 1058 505 1061
rect 622 1061 625 1071
rect 662 1068 673 1071
rect 1110 1068 1118 1071
rect 1166 1068 1174 1071
rect 1182 1068 1201 1071
rect 1206 1068 1222 1071
rect 1302 1068 1321 1071
rect 1438 1068 1449 1071
rect 1542 1068 1550 1071
rect 1582 1068 1590 1071
rect 1606 1068 1625 1071
rect 1822 1068 1838 1071
rect 1846 1068 1857 1071
rect 1974 1068 1982 1071
rect 2018 1068 2030 1071
rect 2326 1071 2329 1078
rect 2318 1068 2329 1071
rect 2342 1071 2345 1081
rect 2846 1078 2857 1081
rect 2966 1078 2974 1081
rect 2846 1072 2849 1078
rect 2342 1068 2350 1071
rect 2642 1068 2649 1071
rect 2670 1068 2678 1071
rect 2822 1068 2841 1071
rect 3014 1068 3033 1071
rect 3038 1068 3062 1071
rect 3078 1068 3105 1071
rect 3174 1068 3182 1071
rect 3222 1068 3241 1071
rect 670 1062 673 1068
rect 974 1062 978 1064
rect 2646 1062 2649 1068
rect 3246 1062 3249 1071
rect 3278 1068 3286 1071
rect 3374 1068 3393 1071
rect 3406 1068 3414 1071
rect 3418 1068 3425 1071
rect 618 1058 625 1061
rect 790 1058 798 1061
rect 1522 1058 1529 1061
rect 1858 1058 1865 1061
rect 2134 1058 2142 1061
rect 2198 1058 2217 1061
rect 2254 1058 2273 1061
rect 2286 1058 2305 1061
rect 2470 1058 2478 1061
rect 2780 1058 2806 1061
rect 2954 1058 2961 1061
rect 3066 1058 3073 1061
rect 3142 1058 3169 1061
rect 3178 1058 3185 1061
rect 3526 1058 3537 1061
rect 262 1048 265 1058
rect 326 1048 329 1058
rect 502 1048 505 1058
rect 542 1048 561 1051
rect 830 1048 849 1051
rect 1218 1048 1225 1051
rect 1286 1048 1294 1051
rect 1642 1048 1646 1052
rect 2286 1048 2289 1058
rect 3526 1057 3530 1058
rect 2574 1048 2585 1051
rect 2610 1048 2617 1051
rect 2938 1048 2942 1052
rect 334 1038 342 1041
rect 414 1038 434 1041
rect 1710 1041 1713 1048
rect 1702 1038 1713 1041
rect 2374 1038 2385 1041
rect 2770 1038 2772 1042
rect 3178 1038 3185 1041
rect 3550 1038 3558 1041
rect 3141 1028 3142 1032
rect 605 1018 606 1022
rect 890 1018 891 1022
rect 954 1018 955 1022
rect 998 1018 1006 1021
rect 1133 1018 1134 1022
rect 1186 1018 1187 1022
rect 1762 1018 1763 1022
rect 2197 1018 2198 1022
rect 2333 1018 2334 1022
rect 2362 1018 2363 1022
rect 2421 1018 2422 1022
rect 2562 1018 2563 1022
rect 480 1003 482 1007
rect 486 1003 489 1007
rect 493 1003 496 1007
rect 1512 1003 1514 1007
rect 1518 1003 1521 1007
rect 1525 1003 1528 1007
rect 2536 1003 2538 1007
rect 2542 1003 2545 1007
rect 2549 1003 2552 1007
rect 749 988 750 992
rect 773 988 774 992
rect 962 988 963 992
rect 1349 988 1350 992
rect 1602 988 1603 992
rect 1781 988 1782 992
rect 1877 988 1878 992
rect 2098 988 2099 992
rect 2850 988 2851 992
rect 3550 988 3558 991
rect 1317 978 1318 982
rect 194 968 201 971
rect 234 968 241 971
rect 78 948 86 951
rect 174 948 182 951
rect 274 948 281 951
rect 330 948 345 951
rect 754 948 769 951
rect 886 951 889 961
rect 870 948 889 951
rect 1006 951 1009 961
rect 1006 948 1041 951
rect 1290 948 1302 951
rect 1486 951 1489 961
rect 2750 958 2761 961
rect 2766 958 2777 961
rect 2774 952 2777 958
rect 1486 948 1505 951
rect 1574 948 1582 951
rect 2282 948 2289 951
rect 2518 948 2534 951
rect 2566 948 2574 951
rect 2642 948 2649 951
rect 2738 948 2753 951
rect 2910 951 2913 961
rect 3414 958 3425 961
rect 2934 951 2937 958
rect 2910 948 2937 951
rect 3030 948 3054 951
rect 54 938 65 941
rect 654 938 665 941
rect 726 941 729 948
rect 718 938 729 941
rect 882 938 889 941
rect 1386 938 1401 941
rect 1586 938 1593 941
rect 1698 938 1705 941
rect 1810 938 1817 941
rect 1926 938 1942 941
rect 2118 941 2121 948
rect 2118 938 2129 941
rect 2198 938 2217 941
rect 2398 938 2406 941
rect 2790 938 2817 941
rect 2830 938 2841 941
rect 2878 938 2889 941
rect 3126 938 3142 941
rect 3190 938 3193 948
rect 3354 938 3361 941
rect 2198 932 2201 938
rect 2186 928 2193 931
rect 2742 928 2745 938
rect 2830 932 2833 938
rect 3510 932 3514 936
rect 13 918 14 922
rect 213 918 214 922
rect 317 918 318 922
rect 1006 918 1022 921
rect 1229 918 1230 922
rect 1901 918 1902 922
rect 2013 918 2014 922
rect 2461 918 2462 922
rect 2692 918 2694 922
rect 992 903 994 907
rect 998 903 1001 907
rect 1005 903 1008 907
rect 2024 903 2026 907
rect 2030 903 2033 907
rect 2037 903 2040 907
rect 3040 903 3042 907
rect 3046 903 3049 907
rect 3053 903 3056 907
rect 413 888 414 892
rect 482 888 497 891
rect 533 888 534 892
rect 733 888 734 892
rect 941 888 942 892
rect 973 888 974 892
rect 1133 888 1134 892
rect 1685 888 1686 892
rect 2845 888 2846 892
rect 3306 888 3308 892
rect 3362 888 3364 892
rect 470 878 478 881
rect 1510 878 1518 881
rect 10 868 17 871
rect 114 868 121 871
rect 166 868 177 871
rect 454 868 462 871
rect 742 868 750 871
rect 982 868 990 871
rect 1006 868 1014 871
rect 1238 868 1254 871
rect 30 858 38 861
rect 54 858 62 861
rect 134 858 153 861
rect 626 858 641 861
rect 678 858 686 861
rect 710 858 718 861
rect 958 858 966 861
rect 1186 858 1201 861
rect 1310 861 1313 871
rect 1334 868 1345 871
rect 1598 871 1601 881
rect 1606 878 1625 881
rect 1970 878 1977 882
rect 2254 878 2265 881
rect 2298 878 2305 881
rect 2406 878 2422 881
rect 2750 878 2761 881
rect 1594 868 1601 871
rect 1622 872 1625 878
rect 1974 872 1977 878
rect 1750 868 1758 871
rect 1306 858 1313 861
rect 1694 861 1697 868
rect 1822 862 1825 871
rect 1642 858 1657 861
rect 1694 858 1713 861
rect 1730 858 1737 861
rect 1854 861 1857 871
rect 1910 868 1918 871
rect 2086 862 2089 871
rect 2734 871 2737 878
rect 2726 868 2737 871
rect 2750 872 2753 878
rect 2766 872 2769 881
rect 2822 878 2830 881
rect 2926 878 2934 882
rect 2998 878 3009 881
rect 3054 878 3070 881
rect 3186 878 3193 881
rect 3198 878 3209 881
rect 2926 872 2929 878
rect 2858 868 2865 871
rect 2886 868 2897 871
rect 3158 871 3161 878
rect 3150 868 3161 871
rect 3218 868 3225 871
rect 3402 868 3409 871
rect 1854 858 1865 861
rect 1942 858 1950 861
rect 2046 858 2054 861
rect 2066 858 2073 861
rect 2226 858 2241 861
rect 2374 858 2382 861
rect 2674 858 2681 861
rect 3178 858 3185 861
rect 3270 858 3286 861
rect 110 848 118 851
rect 134 848 137 858
rect 1162 848 1169 851
rect 1386 848 1390 852
rect 1578 848 1582 852
rect 1822 848 1830 851
rect 2018 848 2033 851
rect 2090 848 2097 851
rect 2106 848 2110 852
rect 2374 848 2377 858
rect 53 838 54 842
rect 86 841 89 848
rect 78 838 89 841
rect 98 838 105 841
rect 122 838 129 841
rect 258 838 265 841
rect 1150 838 1158 841
rect 2330 838 2331 842
rect 3102 838 3113 841
rect 3542 838 3558 841
rect 597 828 598 832
rect 1261 828 1262 832
rect 677 818 678 822
rect 789 818 790 822
rect 818 818 819 822
rect 1074 818 1075 822
rect 1293 818 1294 822
rect 1501 818 1502 822
rect 1714 818 1715 822
rect 1845 818 1846 822
rect 1941 818 1942 822
rect 1997 818 1998 822
rect 2210 818 2211 822
rect 480 803 482 807
rect 486 803 489 807
rect 493 803 496 807
rect 1512 803 1514 807
rect 1518 803 1521 807
rect 1525 803 1528 807
rect 2536 803 2538 807
rect 2542 803 2545 807
rect 2549 803 2552 807
rect 173 788 174 792
rect 397 788 398 792
rect 426 788 427 792
rect 746 788 747 792
rect 1165 788 1166 792
rect 1314 788 1315 792
rect 1510 788 1518 791
rect 1842 788 1843 792
rect 2682 788 2684 792
rect 3066 788 3067 792
rect 3542 788 3550 791
rect 2642 778 2643 782
rect 710 768 721 771
rect 874 768 881 771
rect 1245 768 1246 772
rect 1538 768 1545 771
rect 3181 768 3182 772
rect 718 762 721 768
rect 314 758 318 762
rect 262 751 265 758
rect 262 748 281 751
rect 382 751 385 761
rect 366 748 385 751
rect 438 751 441 761
rect 402 748 425 751
rect 438 748 457 751
rect 530 748 537 751
rect 646 751 649 761
rect 654 758 673 761
rect 630 748 649 751
rect 686 748 702 751
rect 758 751 761 761
rect 758 748 777 751
rect 890 748 902 751
rect 910 748 926 751
rect 1022 751 1025 761
rect 1030 758 1049 761
rect 990 748 1025 751
rect 1134 748 1150 751
rect 1326 748 1334 751
rect 1446 751 1449 761
rect 1490 758 1497 761
rect 1430 748 1449 751
rect 1598 748 1614 751
rect 1918 751 1921 761
rect 2098 758 2105 761
rect 2146 758 2150 762
rect 1902 748 1921 751
rect 2138 748 2145 751
rect 2310 742 2313 751
rect 2486 748 2494 751
rect 2634 748 2641 751
rect 2766 748 2777 751
rect 2790 748 2798 751
rect 2830 751 2833 761
rect 2842 758 2846 762
rect 2814 748 2833 751
rect 2846 748 2854 751
rect 2774 742 2777 748
rect 3058 748 3065 751
rect 3222 748 3230 751
rect 42 738 49 741
rect 254 738 262 741
rect 1174 738 1201 741
rect 1578 738 1585 741
rect 1702 738 1721 741
rect 1890 738 1897 741
rect 2270 738 2278 741
rect 3134 738 3153 741
rect 1522 728 1537 731
rect 1718 728 1721 738
rect 2454 732 2457 738
rect 2190 728 2209 731
rect 2450 728 2457 732
rect 2606 731 2609 738
rect 2606 728 2617 731
rect 3230 728 3233 738
rect 346 718 347 722
rect 478 718 486 721
rect 509 718 510 722
rect 933 718 934 722
rect 957 718 958 722
rect 998 718 1006 721
rect 1114 718 1115 722
rect 1474 718 1476 722
rect 1626 718 1627 722
rect 1645 718 1646 722
rect 992 703 994 707
rect 998 703 1001 707
rect 1005 703 1008 707
rect 2024 703 2026 707
rect 2030 703 2033 707
rect 2037 703 2040 707
rect 3040 703 3042 707
rect 3046 703 3049 707
rect 3053 703 3056 707
rect 162 688 163 692
rect 498 688 505 691
rect 1245 688 1246 692
rect 1941 688 1942 692
rect 3202 688 3204 692
rect 1454 678 1465 681
rect 1506 678 1518 681
rect 202 668 209 671
rect 350 668 358 671
rect 814 668 825 671
rect 910 668 918 671
rect 1758 668 1777 671
rect 1786 668 1809 671
rect 1838 668 1854 671
rect 1894 668 1902 671
rect 2198 671 2201 681
rect 2198 668 2217 671
rect 2854 668 2862 671
rect 3326 668 3334 671
rect 3414 668 3422 671
rect 46 658 65 661
rect 102 658 121 661
rect 286 658 294 661
rect 374 658 393 661
rect 706 658 713 661
rect 774 658 793 661
rect 862 658 881 661
rect 898 658 905 661
rect 922 658 937 661
rect 942 658 958 661
rect 974 658 982 661
rect 1166 658 1185 661
rect 1306 658 1321 661
rect 1338 658 1345 661
rect 1382 658 1390 661
rect 1542 658 1561 661
rect 1794 658 1801 661
rect 1874 658 1881 661
rect 2022 658 2046 661
rect 2474 658 2481 661
rect 2486 658 2505 661
rect 3126 658 3134 661
rect 62 648 65 658
rect 118 648 121 658
rect 390 652 393 658
rect 482 648 505 651
rect 790 648 793 658
rect 862 648 865 658
rect 1166 648 1169 658
rect 1318 648 1321 658
rect 2066 648 2070 652
rect 2430 648 2438 651
rect 285 638 286 642
rect 1218 638 1219 642
rect 1349 638 1350 642
rect 3542 638 3558 641
rect 605 618 606 622
rect 749 618 750 622
rect 805 618 806 622
rect 1154 618 1155 622
rect 1381 618 1382 622
rect 1413 618 1414 622
rect 1988 618 1990 622
rect 2906 618 2907 622
rect 480 603 482 607
rect 486 603 489 607
rect 493 603 496 607
rect 1512 603 1514 607
rect 1518 603 1521 607
rect 1525 603 1528 607
rect 2536 603 2538 607
rect 2542 603 2545 607
rect 2549 603 2552 607
rect 557 588 558 592
rect 818 588 819 592
rect 882 588 883 592
rect 1050 588 1051 592
rect 1210 588 1211 592
rect 1378 588 1379 592
rect 1538 588 1539 592
rect 2621 588 2622 592
rect 2882 588 2883 592
rect 2994 588 2995 592
rect 370 578 371 582
rect 338 568 339 572
rect 733 568 734 572
rect 3086 568 3094 571
rect 262 558 270 561
rect 470 558 489 561
rect 290 548 297 551
rect 462 548 470 551
rect 542 551 545 561
rect 526 548 545 551
rect 558 548 566 551
rect 774 551 777 561
rect 758 548 777 551
rect 830 551 833 561
rect 1082 558 1086 562
rect 798 548 817 551
rect 830 548 849 551
rect 970 548 977 551
rect 982 548 990 551
rect 1086 548 1102 551
rect 1154 548 1161 551
rect 1222 551 1225 561
rect 1346 558 1353 561
rect 2002 558 2006 562
rect 2122 558 2126 562
rect 2274 558 2281 561
rect 1222 548 1241 551
rect 1730 548 1737 551
rect 1766 548 1774 551
rect 1802 548 1817 551
rect 1826 548 1841 551
rect 1942 548 1969 551
rect 2018 548 2041 551
rect 2070 548 2089 551
rect 2146 548 2153 551
rect 54 538 62 541
rect 118 538 126 541
rect 318 541 321 548
rect 798 542 801 548
rect 2382 548 2390 551
rect 2450 548 2457 551
rect 2598 548 2606 551
rect 2714 548 2721 551
rect 2830 548 2849 551
rect 2894 551 2897 561
rect 2894 548 2913 551
rect 3010 548 3025 551
rect 3034 548 3065 551
rect 3174 548 3185 551
rect 3290 548 3297 551
rect 3318 548 3326 551
rect 3366 548 3377 551
rect 3182 542 3185 548
rect 3374 542 3377 548
rect 310 538 321 541
rect 442 538 449 541
rect 570 538 577 541
rect 862 538 870 541
rect 1034 538 1041 541
rect 1254 538 1265 541
rect 1678 538 1686 541
rect 1722 538 1729 541
rect 2498 538 2505 541
rect 2748 538 2750 542
rect 3194 538 3201 541
rect 3318 538 3337 541
rect 582 528 593 531
rect 1774 528 1790 531
rect 2090 528 2097 531
rect 2262 531 2266 533
rect 2262 528 2270 531
rect 2398 531 2402 533
rect 2394 528 2402 531
rect 2530 528 2545 531
rect 3158 528 3166 531
rect 3318 528 3321 538
rect 3346 528 3353 531
rect 2660 518 2662 522
rect 3386 518 3387 522
rect 3550 518 3558 521
rect 992 503 994 507
rect 998 503 1001 507
rect 1005 503 1008 507
rect 2024 503 2026 507
rect 2030 503 2033 507
rect 2037 503 2040 507
rect 3040 503 3042 507
rect 3046 503 3049 507
rect 3053 503 3056 507
rect 418 488 419 492
rect 698 488 699 492
rect 821 488 822 492
rect 2706 488 2713 491
rect 182 478 193 481
rect 302 472 305 481
rect 1822 478 1833 481
rect 154 468 161 471
rect 226 468 233 471
rect 286 468 297 471
rect 370 468 377 471
rect 590 468 598 471
rect 718 468 729 471
rect 198 458 206 461
rect 234 458 241 461
rect 358 458 377 461
rect 538 458 545 461
rect 562 458 577 461
rect 670 458 689 461
rect 730 458 737 461
rect 786 458 793 461
rect 894 461 897 471
rect 966 468 977 471
rect 1134 468 1142 471
rect 1182 468 1190 471
rect 1450 468 1465 471
rect 1510 468 1518 471
rect 1734 468 1745 471
rect 1886 471 1889 481
rect 2206 478 2217 481
rect 2270 478 2281 481
rect 2562 478 2569 481
rect 2870 478 2878 481
rect 1870 468 1889 471
rect 2046 468 2054 471
rect 2458 468 2465 471
rect 2542 468 2577 471
rect 3014 468 3033 471
rect 3142 468 3150 471
rect 3214 468 3233 471
rect 3406 468 3425 471
rect 974 462 977 468
rect 882 458 897 461
rect 994 458 1025 461
rect 1074 458 1081 461
rect 1414 458 1430 461
rect 1702 458 1710 461
rect 2066 458 2073 461
rect 2086 461 2089 468
rect 2086 458 2097 461
rect 2134 458 2142 461
rect 2166 458 2174 461
rect 2294 458 2302 461
rect 2358 458 2374 461
rect 2450 458 2473 461
rect 2590 458 2598 461
rect 2802 458 2817 461
rect 2894 458 2913 461
rect 3046 458 3054 461
rect 3110 458 3118 461
rect 3134 458 3142 461
rect 374 448 377 458
rect 686 452 689 458
rect 2910 452 2913 458
rect 762 448 769 451
rect 1970 448 1974 452
rect 2058 448 2065 451
rect 2130 448 2134 452
rect 3342 448 3353 451
rect 3394 448 3398 452
rect 2165 438 2166 442
rect 1370 418 1374 422
rect 2682 418 2683 422
rect 2850 418 2851 422
rect 480 403 482 407
rect 486 403 489 407
rect 493 403 496 407
rect 1512 403 1514 407
rect 1518 403 1521 407
rect 1525 403 1528 407
rect 2536 403 2538 407
rect 2542 403 2545 407
rect 2549 403 2552 407
rect 210 388 211 392
rect 333 388 334 392
rect 365 388 366 392
rect 413 388 414 392
rect 469 388 470 392
rect 525 388 526 392
rect 610 388 611 392
rect 677 388 678 392
rect 933 388 934 392
rect 965 388 966 392
rect 1130 388 1131 392
rect 1178 388 1179 392
rect 1346 388 1347 392
rect 1642 388 1643 392
rect 1738 388 1739 392
rect 2234 388 2235 392
rect 2594 388 2595 392
rect 2749 388 2750 392
rect 2794 388 2795 392
rect 3146 388 3147 392
rect 3178 388 3179 392
rect 3370 388 3371 392
rect 3506 388 3507 392
rect 1677 368 1678 372
rect 2694 368 2710 371
rect 2858 368 2859 372
rect 558 366 562 368
rect 318 351 321 361
rect 498 358 513 361
rect 546 358 553 361
rect 302 348 321 351
rect 486 348 502 351
rect 558 351 561 361
rect 558 348 577 351
rect 622 351 625 361
rect 622 348 641 351
rect 750 348 758 351
rect 902 348 918 351
rect 1010 348 1017 351
rect 1058 348 1065 351
rect 1202 348 1209 351
rect 1374 351 1377 361
rect 1422 358 1433 361
rect 1370 348 1377 351
rect 1390 348 1398 351
rect 1430 348 1449 351
rect 1654 351 1657 361
rect 3038 358 3046 361
rect 1626 348 1641 351
rect 1654 348 1673 351
rect 1942 351 1945 358
rect 1942 348 1961 351
rect 2034 348 2057 351
rect 2194 348 2201 351
rect 2214 351 2217 358
rect 2214 348 2233 351
rect 2250 348 2257 351
rect 2386 348 2401 351
rect 158 341 161 348
rect 150 338 161 341
rect 290 338 297 341
rect 422 338 433 341
rect 718 338 737 341
rect 1438 338 1446 341
rect 1502 338 1526 341
rect 1622 338 1630 341
rect 1754 338 1761 341
rect 2006 341 2009 348
rect 1990 338 2009 341
rect 2262 338 2289 341
rect 2646 341 2649 351
rect 2766 348 2793 351
rect 2818 348 2825 351
rect 2926 348 2937 351
rect 3170 348 3177 351
rect 3290 348 3297 351
rect 3342 348 3350 351
rect 2934 342 2937 348
rect 2634 338 2649 341
rect 2758 338 2769 341
rect 2914 338 2921 341
rect 3050 338 3070 341
rect 3386 338 3393 341
rect 3454 341 3457 351
rect 3462 348 3470 351
rect 3442 338 3457 341
rect 3462 338 3481 341
rect 3502 338 3529 341
rect 1610 328 1617 331
rect 1622 328 1625 338
rect 2078 332 2081 338
rect 3246 332 3249 338
rect 3318 332 3321 338
rect 2078 328 2086 332
rect 2974 328 2985 331
rect 3242 328 3249 332
rect 3318 328 3326 332
rect 3478 328 3481 338
rect 1261 318 1262 322
rect 1418 318 1419 322
rect 1522 318 1537 321
rect 1580 318 1582 322
rect 992 303 994 307
rect 998 303 1001 307
rect 1005 303 1008 307
rect 2024 303 2026 307
rect 2030 303 2033 307
rect 2037 303 2040 307
rect 3040 303 3042 307
rect 3046 303 3049 307
rect 3053 303 3056 307
rect 178 288 179 292
rect 234 288 235 292
rect 258 288 259 292
rect 445 288 446 292
rect 486 288 494 291
rect 626 288 627 292
rect 1221 288 1222 292
rect 2490 288 2491 292
rect 2754 288 2756 292
rect 3098 288 3099 292
rect 3356 288 3358 292
rect 3509 288 3510 292
rect 966 278 977 281
rect 1070 278 1081 281
rect 1458 278 1465 281
rect 2690 278 2697 281
rect 3038 278 3062 281
rect 3122 278 3129 282
rect 54 268 62 271
rect 150 268 169 271
rect 242 268 249 271
rect 166 262 169 268
rect 34 258 41 261
rect 126 258 134 261
rect 266 258 278 261
rect 290 258 305 261
rect 326 261 329 271
rect 678 268 686 271
rect 726 262 729 271
rect 998 268 1014 271
rect 1042 268 1057 271
rect 1446 268 1454 271
rect 1730 268 1742 271
rect 322 258 329 261
rect 342 258 361 261
rect 486 258 510 261
rect 514 258 521 261
rect 634 258 649 261
rect 686 258 694 261
rect 818 258 825 261
rect 886 258 894 261
rect 918 258 926 261
rect 950 261 953 268
rect 950 258 961 261
rect 1170 258 1185 261
rect 1262 258 1270 261
rect 1286 258 1305 261
rect 1350 258 1361 261
rect 1606 261 1609 268
rect 2142 262 2145 271
rect 2210 268 2217 271
rect 2226 268 2233 271
rect 2318 262 2321 271
rect 2438 271 2441 278
rect 3126 272 3129 278
rect 2438 268 2449 271
rect 2642 268 2649 271
rect 2818 268 2825 271
rect 3082 268 3089 271
rect 3190 271 3193 281
rect 3174 268 3193 271
rect 3270 271 3273 281
rect 3270 268 3297 271
rect 3410 268 3425 271
rect 3478 271 3481 281
rect 3474 268 3481 271
rect 3526 271 3529 281
rect 3534 278 3542 281
rect 3522 268 3529 271
rect 1554 258 1561 261
rect 1590 258 1609 261
rect 1706 258 1721 261
rect 1790 258 1798 261
rect 2034 258 2054 261
rect 2146 258 2172 261
rect 2570 258 2577 261
rect 2590 258 2609 261
rect 2662 261 2665 268
rect 2654 258 2665 261
rect 2670 258 2689 261
rect 2838 258 2865 261
rect 2898 258 2905 261
rect 3238 261 3241 268
rect 3238 258 3249 261
rect 3298 258 3305 261
rect 3454 261 3457 268
rect 3446 258 3457 261
rect 3542 258 3558 261
rect 238 248 246 251
rect 302 248 305 258
rect 310 248 321 251
rect 358 248 361 258
rect 486 248 489 258
rect 686 248 689 258
rect 950 248 961 251
rect 970 248 977 251
rect 1134 248 1142 251
rect 1302 248 1305 258
rect 1350 248 1353 258
rect 1614 248 1625 251
rect 1666 248 1670 252
rect 1790 248 1793 258
rect 2066 248 2070 252
rect 2430 248 2438 251
rect 2590 248 2593 258
rect 2662 248 2673 251
rect 2894 248 2897 258
rect 3126 251 3129 258
rect 3126 248 3137 251
rect 3166 251 3169 258
rect 3158 248 3169 251
rect 3446 248 3457 251
rect 318 242 321 248
rect 1350 242 1354 244
rect 741 238 742 242
rect 2214 238 2222 241
rect 3490 238 3491 242
rect 2030 228 2038 231
rect 1317 218 1318 222
rect 1538 218 1539 222
rect 1637 218 1638 222
rect 3306 218 3307 222
rect 3346 218 3348 222
rect 480 203 482 207
rect 486 203 489 207
rect 493 203 496 207
rect 1512 203 1514 207
rect 1518 203 1521 207
rect 1525 203 1528 207
rect 2536 203 2538 207
rect 2542 203 2545 207
rect 2549 203 2552 207
rect 362 188 363 192
rect 509 188 510 192
rect 613 188 614 192
rect 917 188 918 192
rect 1026 188 1030 192
rect 1074 188 1075 192
rect 1605 188 1606 192
rect 1629 188 1630 192
rect 1661 188 1662 192
rect 1834 188 1835 192
rect 1866 188 1867 192
rect 2277 188 2278 192
rect 2338 188 2339 192
rect 2469 188 2470 192
rect 2510 188 2518 191
rect 2564 188 2566 192
rect 2698 188 2700 192
rect 2773 188 2774 192
rect 2890 188 2891 192
rect 3413 188 3414 192
rect 1458 178 1459 182
rect 298 168 305 171
rect 570 168 571 172
rect 758 168 766 171
rect 861 168 862 172
rect 1214 168 1225 171
rect 2350 168 2374 171
rect 3186 168 3187 172
rect 1214 162 1217 168
rect 654 158 673 161
rect 126 148 134 151
rect 226 148 233 151
rect 258 148 265 151
rect 342 148 358 151
rect 634 148 641 151
rect 710 151 713 161
rect 974 158 982 161
rect 1222 158 1233 161
rect 1414 158 1425 161
rect 1582 158 1593 161
rect 1902 158 1918 161
rect 2438 161 2441 168
rect 2430 158 2441 161
rect 2622 158 2633 161
rect 3034 158 3038 162
rect 3162 158 3169 161
rect 3390 158 3401 161
rect 694 148 713 151
rect 918 148 945 151
rect 1402 148 1417 151
rect 1554 148 1561 151
rect 1614 148 1625 151
rect 1758 148 1766 151
rect 2014 148 2038 151
rect 2198 148 2214 151
rect 2254 148 2262 151
rect 2318 148 2329 151
rect 2454 151 2457 158
rect 2502 151 2505 158
rect 2454 148 2465 151
rect 2494 148 2505 151
rect 2606 148 2625 151
rect 2638 148 2657 151
rect 2850 148 2857 151
rect 3014 148 3022 151
rect 3058 148 3097 151
rect 3342 148 3353 151
rect 3414 148 3422 151
rect 3446 148 3462 151
rect 3502 148 3521 151
rect 22 138 30 141
rect 86 138 94 141
rect 342 141 345 148
rect 1614 142 1617 148
rect 290 138 297 141
rect 334 138 345 141
rect 1194 138 1201 141
rect 1258 138 1265 141
rect 1366 138 1382 141
rect 1494 138 1502 141
rect 1550 138 1566 141
rect 1718 138 1737 141
rect 1946 138 1953 141
rect 2094 138 2113 141
rect 2222 141 2225 148
rect 2222 138 2241 141
rect 2326 138 2329 148
rect 2582 138 2590 141
rect 2654 138 2657 148
rect 2674 138 2681 141
rect 2742 138 2750 141
rect 3006 138 3014 141
rect 3094 138 3097 148
rect 3342 142 3345 148
rect 3118 138 3137 141
rect 3238 138 3257 141
rect 3270 138 3305 141
rect 3458 138 3473 141
rect 3490 138 3497 141
rect 1390 128 1398 131
rect 1502 128 1510 131
rect 3270 128 3273 138
rect 1980 118 1982 122
rect 3338 118 3339 122
rect 992 103 994 107
rect 998 103 1001 107
rect 1005 103 1008 107
rect 2024 103 2026 107
rect 2030 103 2033 107
rect 2037 103 2040 107
rect 3040 103 3042 107
rect 3046 103 3049 107
rect 3053 103 3056 107
rect 354 88 355 92
rect 426 88 427 92
rect 478 88 494 91
rect 778 88 779 92
rect 858 88 859 92
rect 890 88 891 92
rect 1156 88 1158 92
rect 1596 88 1598 92
rect 2092 88 2094 92
rect 2188 88 2190 92
rect 2508 88 2510 92
rect 2892 88 2894 92
rect 3098 88 3100 92
rect 3221 88 3222 92
rect 3268 88 3270 92
rect 1002 78 1009 81
rect 22 68 33 71
rect 434 68 441 71
rect 490 68 513 71
rect 934 71 937 78
rect 842 68 849 71
rect 926 68 937 71
rect 1670 71 1673 81
rect 1686 78 1697 81
rect 1694 72 1697 78
rect 1670 68 1689 71
rect 1734 71 1737 81
rect 1794 78 1809 81
rect 2026 78 2033 81
rect 1734 68 1753 71
rect 1998 68 2030 71
rect 30 62 33 68
rect 2158 62 2161 71
rect 2214 71 2217 81
rect 2278 78 2286 81
rect 3054 78 3062 81
rect 3138 78 3145 81
rect 2210 68 2217 71
rect 2410 68 2425 71
rect 2430 68 2438 71
rect 2470 68 2478 71
rect 2566 71 2569 78
rect 2554 68 2561 71
rect 2566 68 2577 71
rect 2730 68 2737 71
rect 2778 68 2793 71
rect 2802 68 2809 71
rect 3038 71 3041 78
rect 3038 68 3049 71
rect 3206 68 3214 71
rect 3366 68 3374 71
rect 274 58 281 61
rect 686 58 705 61
rect 730 58 737 61
rect 974 58 1009 61
rect 1046 58 1065 61
rect 1090 58 1097 61
rect 1190 58 1201 61
rect 1206 58 1222 61
rect 1274 58 1281 61
rect 1324 58 1326 62
rect 1390 58 1414 61
rect 1422 58 1430 61
rect 1502 58 1518 61
rect 1630 58 1649 61
rect 1694 58 1721 61
rect 1750 58 1761 61
rect 1790 58 1798 61
rect 2350 58 2358 61
rect 2434 58 2441 61
rect 2462 58 2470 61
rect 2582 58 2598 61
rect 2942 58 2950 61
rect 3006 58 3041 61
rect 574 48 593 51
rect 702 48 705 58
rect 1006 48 1009 58
rect 1062 48 1065 58
rect 1258 48 1262 52
rect 1798 48 1806 51
rect 1886 48 1897 51
rect 2350 48 2353 58
rect 2626 48 2633 51
rect 1077 38 1078 42
rect 1830 38 1838 41
rect 2836 38 2838 42
rect 2965 38 2966 42
rect 717 28 718 32
rect 2365 28 2366 32
rect 2610 28 2611 32
rect 480 3 482 7
rect 486 3 489 7
rect 493 3 496 7
rect 1512 3 1514 7
rect 1518 3 1521 7
rect 1525 3 1528 7
rect 2536 3 2538 7
rect 2542 3 2545 7
rect 2549 3 2552 7
<< m2contact >>
rect 994 3303 998 3307
rect 1001 3303 1005 3307
rect 2026 3303 2030 3307
rect 2033 3303 2037 3307
rect 3042 3303 3046 3307
rect 3049 3303 3053 3307
rect 182 3288 186 3292
rect 326 3288 330 3292
rect 414 3288 418 3292
rect 502 3288 506 3292
rect 534 3288 538 3292
rect 926 3288 930 3292
rect 1350 3288 1354 3292
rect 1630 3288 1634 3292
rect 2014 3288 2018 3292
rect 2054 3288 2058 3292
rect 2102 3288 2106 3292
rect 2126 3288 2130 3292
rect 2174 3288 2178 3292
rect 2278 3288 2282 3292
rect 2302 3288 2306 3292
rect 2326 3288 2330 3292
rect 2350 3288 2354 3292
rect 2390 3288 2394 3292
rect 2406 3288 2410 3292
rect 2430 3288 2434 3292
rect 2470 3288 2474 3292
rect 2494 3288 2498 3292
rect 2558 3288 2562 3292
rect 2582 3288 2586 3292
rect 2606 3288 2610 3292
rect 2630 3288 2634 3292
rect 2686 3288 2690 3292
rect 2950 3288 2954 3292
rect 2974 3288 2978 3292
rect 2998 3288 3002 3292
rect 3022 3288 3026 3292
rect 3062 3288 3066 3292
rect 3126 3288 3130 3292
rect 3150 3288 3154 3292
rect 3190 3288 3194 3292
rect 3214 3288 3218 3292
rect 3238 3288 3242 3292
rect 3318 3288 3322 3292
rect 3342 3288 3346 3292
rect 174 3278 178 3282
rect 222 3278 226 3282
rect 390 3278 394 3282
rect 470 3278 474 3282
rect 654 3278 658 3282
rect 110 3268 114 3272
rect 134 3268 138 3272
rect 254 3268 258 3272
rect 462 3268 466 3272
rect 622 3268 626 3272
rect 774 3278 778 3282
rect 782 3278 786 3282
rect 886 3278 890 3282
rect 894 3278 898 3282
rect 958 3278 962 3282
rect 998 3278 1002 3282
rect 1014 3278 1018 3282
rect 678 3268 682 3272
rect 694 3268 698 3272
rect 766 3268 770 3272
rect 854 3268 858 3272
rect 870 3268 874 3272
rect 886 3268 890 3272
rect 910 3268 914 3272
rect 958 3268 962 3272
rect 1006 3268 1010 3272
rect 1038 3268 1042 3272
rect 1078 3268 1082 3272
rect 1094 3268 1098 3272
rect 1118 3278 1122 3282
rect 1174 3278 1178 3282
rect 1382 3278 1386 3282
rect 1462 3278 1466 3282
rect 1654 3278 1658 3282
rect 1686 3278 1690 3282
rect 1806 3278 1810 3282
rect 1342 3268 1346 3272
rect 1454 3268 1458 3272
rect 1478 3268 1482 3272
rect 1518 3268 1522 3272
rect 1566 3268 1570 3272
rect 1646 3268 1650 3272
rect 1702 3268 1706 3272
rect 2078 3278 2082 3282
rect 2150 3278 2154 3282
rect 2182 3278 2186 3282
rect 2238 3278 2242 3282
rect 2374 3278 2378 3282
rect 2518 3278 2522 3282
rect 2662 3278 2666 3282
rect 2694 3278 2698 3282
rect 3070 3278 3074 3282
rect 3110 3278 3114 3282
rect 3382 3278 3386 3282
rect 3510 3278 3514 3282
rect 1830 3268 1834 3272
rect 1846 3268 1850 3272
rect 1902 3268 1906 3272
rect 1918 3268 1922 3272
rect 1934 3268 1938 3272
rect 2078 3268 2082 3272
rect 2110 3268 2114 3272
rect 2126 3268 2130 3272
rect 2502 3268 2506 3272
rect 2638 3268 2642 3272
rect 2654 3268 2658 3272
rect 2782 3268 2786 3272
rect 2814 3268 2818 3272
rect 2854 3268 2858 3272
rect 2894 3268 2898 3272
rect 3310 3268 3314 3272
rect 3382 3268 3386 3272
rect 3438 3268 3442 3272
rect 3462 3268 3466 3272
rect 3486 3268 3490 3272
rect 3518 3268 3522 3272
rect 94 3259 98 3263
rect 126 3258 130 3262
rect 142 3258 146 3262
rect 158 3258 162 3262
rect 198 3258 202 3262
rect 206 3258 210 3262
rect 262 3258 266 3262
rect 342 3258 346 3262
rect 366 3258 370 3262
rect 398 3258 402 3262
rect 422 3258 426 3262
rect 478 3258 482 3262
rect 518 3258 522 3262
rect 606 3259 610 3263
rect 638 3258 642 3262
rect 662 3258 666 3262
rect 686 3258 690 3262
rect 702 3258 706 3262
rect 734 3258 738 3262
rect 742 3258 746 3262
rect 758 3258 762 3262
rect 790 3258 794 3262
rect 862 3258 866 3262
rect 902 3258 906 3262
rect 918 3258 922 3262
rect 942 3258 946 3262
rect 974 3258 978 3262
rect 1046 3258 1050 3262
rect 1070 3258 1074 3262
rect 1086 3258 1090 3262
rect 1110 3258 1114 3262
rect 1198 3258 1202 3262
rect 1270 3258 1274 3262
rect 1294 3258 1298 3262
rect 1334 3258 1338 3262
rect 1366 3258 1370 3262
rect 1470 3258 1474 3262
rect 1486 3258 1490 3262
rect 1510 3258 1514 3262
rect 1590 3258 1594 3262
rect 1638 3258 1642 3262
rect 1670 3258 1674 3262
rect 1726 3258 1730 3262
rect 1790 3258 1794 3262
rect 1814 3258 1818 3262
rect 1838 3258 1842 3262
rect 1854 3258 1858 3262
rect 1950 3259 1954 3263
rect 2038 3258 2042 3262
rect 2062 3258 2066 3262
rect 2086 3258 2090 3262
rect 2134 3258 2138 3262
rect 2158 3258 2162 3262
rect 2198 3258 2202 3262
rect 2214 3258 2218 3262
rect 2254 3258 2258 3262
rect 2262 3258 2266 3262
rect 2286 3258 2290 3262
rect 2310 3258 2314 3262
rect 2334 3258 2338 3262
rect 2358 3258 2362 3262
rect 2422 3258 2426 3262
rect 2446 3258 2450 3262
rect 2454 3258 2458 3262
rect 2478 3258 2482 3262
rect 2502 3258 2506 3262
rect 2526 3258 2530 3262
rect 2558 3258 2562 3262
rect 2590 3258 2594 3262
rect 2614 3258 2618 3262
rect 2670 3258 2674 3262
rect 2694 3258 2698 3262
rect 2710 3258 2714 3262
rect 2774 3258 2778 3262
rect 2830 3258 2834 3262
rect 2846 3258 2850 3262
rect 2886 3259 2890 3263
rect 2958 3258 2962 3262
rect 2982 3258 2986 3262
rect 3006 3258 3010 3262
rect 3030 3258 3034 3262
rect 3086 3258 3090 3262
rect 3094 3258 3098 3262
rect 3110 3258 3114 3262
rect 3126 3258 3130 3262
rect 3166 3258 3170 3262
rect 3174 3258 3178 3262
rect 3198 3258 3202 3262
rect 3222 3258 3226 3262
rect 3246 3258 3250 3262
rect 3334 3258 3338 3262
rect 3358 3258 3362 3262
rect 3366 3258 3370 3262
rect 3382 3258 3386 3262
rect 3398 3258 3402 3262
rect 3494 3258 3498 3262
rect 3510 3258 3514 3262
rect 3526 3258 3530 3262
rect 214 3248 218 3252
rect 350 3248 354 3252
rect 358 3248 362 3252
rect 430 3248 434 3252
rect 726 3248 730 3252
rect 926 3248 930 3252
rect 1054 3248 1058 3252
rect 1494 3248 1498 3252
rect 1510 3248 1514 3252
rect 1870 3248 1874 3252
rect 1894 3248 1898 3252
rect 2126 3248 2130 3252
rect 6 3238 10 3242
rect 30 3238 34 3242
rect 542 3238 546 3242
rect 558 3238 562 3242
rect 1022 3238 1026 3242
rect 1070 3238 1074 3242
rect 1326 3238 1330 3242
rect 1398 3238 1402 3242
rect 1766 3238 1770 3242
rect 2230 3248 2234 3252
rect 2398 3248 2402 3252
rect 2830 3248 2834 3252
rect 2846 3248 2850 3252
rect 3118 3248 3122 3252
rect 3414 3248 3418 3252
rect 3422 3248 3426 3252
rect 3446 3248 3450 3252
rect 3470 3248 3474 3252
rect 2222 3238 2226 3242
rect 2718 3238 2722 3242
rect 3086 3238 3090 3242
rect 3134 3238 3138 3242
rect 2246 3228 2250 3232
rect 3398 3228 3402 3232
rect 318 3218 322 3222
rect 718 3218 722 3222
rect 966 3218 970 3222
rect 3430 3218 3434 3222
rect 3454 3218 3458 3222
rect 3478 3218 3482 3222
rect 3542 3218 3546 3222
rect 482 3203 486 3207
rect 489 3203 493 3207
rect 1514 3203 1518 3207
rect 1521 3203 1525 3207
rect 2538 3203 2542 3207
rect 2545 3203 2549 3207
rect 102 3188 106 3192
rect 174 3188 178 3192
rect 334 3188 338 3192
rect 366 3188 370 3192
rect 910 3188 914 3192
rect 934 3188 938 3192
rect 974 3188 978 3192
rect 1110 3188 1114 3192
rect 1262 3188 1266 3192
rect 1574 3188 1578 3192
rect 1838 3188 1842 3192
rect 2438 3188 2442 3192
rect 2638 3188 2642 3192
rect 2718 3188 2722 3192
rect 2774 3188 2778 3192
rect 2934 3188 2938 3192
rect 3294 3188 3298 3192
rect 1966 3178 1970 3182
rect 2974 3178 2978 3182
rect 3206 3178 3210 3182
rect 94 3168 98 3172
rect 710 3168 714 3172
rect 814 3168 818 3172
rect 1206 3168 1210 3172
rect 1254 3168 1258 3172
rect 1406 3168 1410 3172
rect 1782 3168 1786 3172
rect 2110 3168 2114 3172
rect 2670 3168 2674 3172
rect 30 3158 34 3162
rect 14 3148 18 3152
rect 38 3148 42 3152
rect 78 3158 82 3162
rect 110 3158 114 3162
rect 566 3158 570 3162
rect 582 3158 586 3162
rect 598 3158 602 3162
rect 638 3158 642 3162
rect 670 3158 674 3162
rect 798 3158 802 3162
rect 830 3158 834 3162
rect 878 3158 882 3162
rect 918 3158 922 3162
rect 950 3158 954 3162
rect 1182 3158 1186 3162
rect 1190 3158 1194 3162
rect 1238 3158 1242 3162
rect 1286 3158 1290 3162
rect 1310 3158 1314 3162
rect 1734 3158 1738 3162
rect 1822 3158 1826 3162
rect 2270 3158 2274 3162
rect 2342 3158 2346 3162
rect 2478 3158 2482 3162
rect 2494 3158 2498 3162
rect 2702 3158 2706 3162
rect 2710 3158 2714 3162
rect 3054 3158 3058 3162
rect 3222 3158 3226 3162
rect 3278 3158 3282 3162
rect 3310 3158 3314 3162
rect 102 3148 106 3152
rect 150 3148 154 3152
rect 182 3148 186 3152
rect 254 3148 258 3152
rect 278 3147 282 3151
rect 310 3148 314 3152
rect 342 3148 346 3152
rect 406 3148 410 3152
rect 494 3148 498 3152
rect 550 3148 554 3152
rect 582 3148 586 3152
rect 606 3148 610 3152
rect 630 3148 634 3152
rect 678 3148 682 3152
rect 742 3148 746 3152
rect 766 3148 770 3152
rect 798 3148 802 3152
rect 814 3148 818 3152
rect 838 3148 842 3152
rect 974 3148 978 3152
rect 6 3138 10 3142
rect 30 3138 34 3142
rect 78 3138 82 3142
rect 134 3138 138 3142
rect 158 3138 162 3142
rect 174 3138 178 3142
rect 206 3138 210 3142
rect 294 3138 298 3142
rect 318 3138 322 3142
rect 406 3138 410 3142
rect 446 3138 450 3142
rect 518 3138 522 3142
rect 542 3138 546 3142
rect 574 3138 578 3142
rect 654 3138 658 3142
rect 734 3138 738 3142
rect 774 3138 778 3142
rect 1038 3147 1042 3151
rect 1118 3148 1122 3152
rect 1166 3148 1170 3152
rect 1190 3148 1194 3152
rect 1246 3148 1250 3152
rect 1278 3148 1282 3152
rect 1350 3148 1354 3152
rect 1374 3148 1378 3152
rect 1430 3148 1434 3152
rect 1518 3148 1522 3152
rect 1662 3148 1666 3152
rect 1686 3148 1690 3152
rect 1702 3148 1706 3152
rect 1718 3148 1722 3152
rect 1742 3148 1746 3152
rect 1758 3148 1762 3152
rect 1838 3148 1842 3152
rect 1846 3148 1850 3152
rect 1870 3148 1874 3152
rect 806 3138 810 3142
rect 862 3138 866 3142
rect 894 3138 898 3142
rect 942 3138 946 3142
rect 966 3138 970 3142
rect 1022 3138 1026 3142
rect 1134 3138 1138 3142
rect 1158 3138 1162 3142
rect 1214 3138 1218 3142
rect 1270 3138 1274 3142
rect 1294 3138 1298 3142
rect 1342 3138 1346 3142
rect 1382 3138 1386 3142
rect 1438 3138 1442 3142
rect 1510 3138 1514 3142
rect 1606 3138 1610 3142
rect 1654 3138 1658 3142
rect 1694 3138 1698 3142
rect 1902 3147 1906 3151
rect 1934 3148 1938 3152
rect 1974 3148 1978 3152
rect 2006 3148 2010 3152
rect 2046 3147 2050 3151
rect 2134 3148 2138 3152
rect 2142 3148 2146 3152
rect 2222 3148 2226 3152
rect 2246 3148 2250 3152
rect 2294 3148 2298 3152
rect 2326 3148 2330 3152
rect 2342 3148 2346 3152
rect 1742 3138 1746 3142
rect 1782 3138 1786 3142
rect 1806 3140 1810 3144
rect 1814 3138 1818 3142
rect 1846 3138 1850 3142
rect 1982 3138 1986 3142
rect 2030 3138 2034 3142
rect 2166 3138 2170 3142
rect 2190 3138 2194 3142
rect 2254 3138 2258 3142
rect 2270 3138 2274 3142
rect 2310 3138 2314 3142
rect 2374 3147 2378 3151
rect 2486 3148 2490 3152
rect 2526 3148 2530 3152
rect 2574 3147 2578 3151
rect 2646 3148 2650 3152
rect 2686 3148 2690 3152
rect 2734 3148 2738 3152
rect 2750 3148 2754 3152
rect 2782 3148 2786 3152
rect 2798 3148 2802 3152
rect 2830 3148 2834 3152
rect 2862 3147 2866 3151
rect 2894 3148 2898 3152
rect 2958 3148 2962 3152
rect 2974 3148 2978 3152
rect 3006 3147 3010 3151
rect 3038 3148 3042 3152
rect 3110 3148 3114 3152
rect 3142 3147 3146 3151
rect 3174 3148 3178 3152
rect 3254 3148 3258 3152
rect 3334 3148 3338 3152
rect 3358 3148 3362 3152
rect 3382 3148 3386 3152
rect 3438 3148 3442 3152
rect 3462 3148 3466 3152
rect 3526 3148 3530 3152
rect 3534 3148 3538 3152
rect 2358 3138 2362 3142
rect 2390 3138 2394 3142
rect 2582 3138 2586 3142
rect 2654 3138 2658 3142
rect 2678 3138 2682 3142
rect 2790 3138 2794 3142
rect 3078 3138 3082 3142
rect 3126 3138 3130 3142
rect 3326 3138 3330 3142
rect 3398 3138 3402 3142
rect 3502 3138 3506 3142
rect 3558 3138 3562 3142
rect 54 3128 58 3132
rect 118 3128 122 3132
rect 142 3128 146 3132
rect 174 3128 178 3132
rect 206 3128 210 3132
rect 358 3128 362 3132
rect 462 3128 466 3132
rect 502 3128 506 3132
rect 606 3128 610 3132
rect 622 3128 626 3132
rect 678 3128 682 3132
rect 694 3128 698 3132
rect 718 3128 722 3132
rect 750 3128 754 3132
rect 766 3128 770 3132
rect 854 3128 858 3132
rect 910 3128 914 3132
rect 990 3128 994 3132
rect 1118 3128 1122 3132
rect 1150 3128 1154 3132
rect 1230 3128 1234 3132
rect 1350 3128 1354 3132
rect 1366 3128 1370 3132
rect 1398 3128 1402 3132
rect 1406 3128 1410 3132
rect 1462 3128 1466 3132
rect 1598 3128 1602 3132
rect 1662 3128 1666 3132
rect 1678 3128 1682 3132
rect 1742 3128 1746 3132
rect 1758 3128 1762 3132
rect 1854 3128 1858 3132
rect 1998 3128 2002 3132
rect 2118 3128 2122 3132
rect 2134 3128 2138 3132
rect 2174 3128 2178 3132
rect 2206 3128 2210 3132
rect 2230 3128 2234 3132
rect 2462 3128 2466 3132
rect 2470 3128 2474 3132
rect 2494 3128 2498 3132
rect 2510 3128 2514 3132
rect 2670 3128 2674 3132
rect 2702 3128 2706 3132
rect 2750 3128 2754 3132
rect 2814 3128 2818 3132
rect 2958 3128 2962 3132
rect 3094 3128 3098 3132
rect 3230 3128 3234 3132
rect 3238 3128 3242 3132
rect 3350 3128 3354 3132
rect 3358 3128 3362 3132
rect 3374 3128 3378 3132
rect 214 3118 218 3122
rect 366 3118 370 3122
rect 470 3118 474 3122
rect 566 3118 570 3122
rect 670 3118 674 3122
rect 726 3118 730 3122
rect 846 3118 850 3122
rect 950 3118 954 3122
rect 1102 3118 1106 3122
rect 1142 3118 1146 3122
rect 1590 3118 1594 3122
rect 1638 3118 1642 3122
rect 2182 3118 2186 3122
rect 2238 3118 2242 3122
rect 2262 3118 2266 3122
rect 2302 3118 2306 3122
rect 2454 3118 2458 3122
rect 2518 3118 2522 3122
rect 2926 3118 2930 3122
rect 3078 3118 3082 3122
rect 3342 3118 3346 3122
rect 3390 3118 3394 3122
rect 994 3103 998 3107
rect 1001 3103 1005 3107
rect 2026 3103 2030 3107
rect 2033 3103 2037 3107
rect 3042 3103 3046 3107
rect 3049 3103 3053 3107
rect 46 3088 50 3092
rect 134 3088 138 3092
rect 166 3088 170 3092
rect 294 3088 298 3092
rect 350 3088 354 3092
rect 398 3088 402 3092
rect 494 3088 498 3092
rect 606 3088 610 3092
rect 822 3088 826 3092
rect 902 3088 906 3092
rect 1062 3088 1066 3092
rect 1206 3088 1210 3092
rect 1230 3088 1234 3092
rect 1406 3088 1410 3092
rect 1462 3088 1466 3092
rect 1494 3088 1498 3092
rect 1574 3088 1578 3092
rect 1646 3088 1650 3092
rect 1670 3088 1674 3092
rect 1814 3088 1818 3092
rect 1878 3088 1882 3092
rect 1958 3088 1962 3092
rect 1998 3088 2002 3092
rect 2134 3088 2138 3092
rect 2294 3088 2298 3092
rect 2422 3088 2426 3092
rect 2534 3088 2538 3092
rect 2590 3088 2594 3092
rect 2686 3088 2690 3092
rect 2798 3088 2802 3092
rect 2838 3088 2842 3092
rect 3014 3088 3018 3092
rect 3182 3088 3186 3092
rect 3310 3088 3314 3092
rect 3382 3088 3386 3092
rect 3510 3088 3514 3092
rect 3550 3088 3554 3092
rect 6 3078 10 3082
rect 22 3078 26 3082
rect 30 3068 34 3072
rect 54 3068 58 3072
rect 70 3068 74 3072
rect 86 3078 90 3082
rect 238 3078 242 3082
rect 326 3078 330 3082
rect 358 3078 362 3082
rect 382 3078 386 3082
rect 142 3068 146 3072
rect 174 3068 178 3072
rect 198 3068 202 3072
rect 222 3068 226 3072
rect 246 3068 250 3072
rect 286 3068 290 3072
rect 342 3068 346 3072
rect 478 3078 482 3082
rect 598 3078 602 3082
rect 718 3078 722 3082
rect 734 3078 738 3082
rect 814 3078 818 3082
rect 862 3078 866 3082
rect 870 3078 874 3082
rect 910 3078 914 3082
rect 926 3078 930 3082
rect 958 3078 962 3082
rect 1150 3078 1154 3082
rect 1158 3078 1162 3082
rect 1214 3078 1218 3082
rect 1222 3078 1226 3082
rect 1254 3078 1258 3082
rect 1350 3078 1354 3082
rect 1390 3078 1394 3082
rect 1398 3078 1402 3082
rect 1446 3078 1450 3082
rect 1502 3078 1506 3082
rect 1542 3078 1546 3082
rect 1566 3078 1570 3082
rect 1582 3078 1586 3082
rect 1614 3078 1618 3082
rect 1678 3078 1682 3082
rect 1710 3078 1714 3082
rect 1822 3078 1826 3082
rect 1886 3078 1890 3082
rect 2006 3078 2010 3082
rect 2046 3078 2050 3082
rect 462 3068 466 3072
rect 558 3068 562 3072
rect 614 3068 618 3072
rect 646 3068 650 3072
rect 678 3068 682 3072
rect 686 3068 690 3072
rect 830 3068 834 3072
rect 934 3068 938 3072
rect 966 3068 970 3072
rect 1038 3068 1042 3072
rect 1046 3068 1050 3072
rect 1070 3068 1074 3072
rect 1078 3068 1082 3072
rect 1102 3068 1106 3072
rect 1134 3068 1138 3072
rect 1150 3068 1154 3072
rect 1238 3068 1242 3072
rect 1286 3068 1290 3072
rect 1326 3068 1330 3072
rect 1342 3068 1346 3072
rect 1414 3068 1418 3072
rect 1470 3068 1474 3072
rect 1486 3068 1490 3072
rect 1582 3068 1586 3072
rect 1622 3068 1626 3072
rect 1662 3068 1666 3072
rect 1694 3068 1698 3072
rect 1702 3068 1706 3072
rect 1758 3068 1762 3072
rect 1806 3068 1810 3072
rect 1830 3068 1834 3072
rect 1846 3068 1850 3072
rect 1886 3068 1890 3072
rect 1926 3068 1930 3072
rect 1974 3068 1978 3072
rect 1990 3068 1994 3072
rect 2014 3068 2018 3072
rect 2062 3078 2066 3082
rect 2086 3078 2090 3082
rect 2142 3078 2146 3082
rect 2150 3078 2154 3082
rect 2230 3078 2234 3082
rect 2358 3078 2362 3082
rect 2438 3078 2442 3082
rect 2510 3078 2514 3082
rect 2542 3078 2546 3082
rect 2070 3068 2074 3072
rect 2094 3068 2098 3072
rect 2102 3068 2106 3072
rect 2126 3068 2130 3072
rect 2158 3068 2162 3072
rect 2190 3068 2194 3072
rect 2262 3068 2266 3072
rect 2270 3068 2274 3072
rect 2374 3068 2378 3072
rect 2390 3068 2394 3072
rect 2446 3068 2450 3072
rect 2454 3068 2458 3072
rect 2470 3068 2474 3072
rect 2494 3068 2498 3072
rect 2526 3068 2530 3072
rect 2566 3068 2570 3072
rect 2702 3068 2706 3072
rect 2830 3068 2834 3072
rect 2854 3078 2858 3082
rect 2974 3078 2978 3082
rect 2990 3078 2994 3082
rect 3022 3078 3026 3082
rect 3062 3078 3066 3082
rect 3086 3078 3090 3082
rect 3214 3078 3218 3082
rect 3246 3078 3250 3082
rect 3318 3078 3322 3082
rect 3390 3078 3394 3082
rect 3526 3078 3530 3082
rect 2886 3068 2890 3072
rect 3006 3068 3010 3072
rect 3030 3068 3034 3072
rect 3070 3068 3074 3072
rect 3126 3068 3130 3072
rect 3198 3068 3202 3072
rect 3214 3068 3218 3072
rect 3334 3068 3338 3072
rect 3366 3068 3370 3072
rect 3422 3068 3426 3072
rect 3438 3068 3442 3072
rect 22 3058 26 3062
rect 62 3058 66 3062
rect 102 3058 106 3062
rect 118 3058 122 3062
rect 150 3058 154 3062
rect 214 3058 218 3062
rect 254 3058 258 3062
rect 310 3058 314 3062
rect 334 3058 338 3062
rect 366 3058 370 3062
rect 414 3058 418 3062
rect 438 3058 442 3062
rect 454 3058 458 3062
rect 470 3058 474 3062
rect 566 3059 570 3063
rect 622 3058 626 3062
rect 670 3058 674 3062
rect 694 3058 698 3062
rect 750 3058 754 3062
rect 798 3058 802 3062
rect 838 3058 842 3062
rect 846 3058 850 3062
rect 886 3058 890 3062
rect 942 3058 946 3062
rect 958 3058 962 3062
rect 1030 3058 1034 3062
rect 1054 3058 1058 3062
rect 1126 3058 1130 3062
rect 1150 3058 1154 3062
rect 1190 3058 1194 3062
rect 1246 3058 1250 3062
rect 1270 3058 1274 3062
rect 1310 3058 1314 3062
rect 1366 3058 1370 3062
rect 1374 3058 1378 3062
rect 1422 3058 1426 3062
rect 1430 3058 1434 3062
rect 1478 3058 1482 3062
rect 1526 3058 1530 3062
rect 1630 3058 1634 3062
rect 1654 3058 1658 3062
rect 1726 3058 1730 3062
rect 1790 3058 1794 3062
rect 1798 3058 1802 3062
rect 1902 3058 1906 3062
rect 1926 3058 1930 3062
rect 1982 3058 1986 3062
rect 2014 3058 2018 3062
rect 2078 3058 2082 3062
rect 2110 3058 2114 3062
rect 2118 3058 2122 3062
rect 2198 3058 2202 3062
rect 2214 3058 2218 3062
rect 2286 3058 2290 3062
rect 2350 3058 2354 3062
rect 2406 3058 2410 3062
rect 2454 3058 2458 3062
rect 2486 3058 2490 3062
rect 2502 3058 2506 3062
rect 2518 3058 2522 3062
rect 2574 3058 2578 3062
rect 2630 3058 2634 3062
rect 2654 3058 2658 3062
rect 2718 3059 2722 3063
rect 2750 3058 2754 3062
rect 2814 3058 2818 3062
rect 2822 3058 2826 3062
rect 2870 3058 2874 3062
rect 2910 3058 2914 3062
rect 2998 3058 3002 3062
rect 3038 3058 3042 3062
rect 3118 3059 3122 3063
rect 3190 3058 3194 3062
rect 3246 3059 3250 3063
rect 3438 3058 3442 3062
rect 3534 3058 3538 3062
rect 190 3048 194 3052
rect 270 3048 274 3052
rect 422 3048 426 3052
rect 630 3048 634 3052
rect 774 3048 778 3052
rect 782 3048 786 3052
rect 798 3048 802 3052
rect 918 3048 922 3052
rect 1086 3048 1090 3052
rect 1094 3048 1098 3052
rect 1118 3048 1122 3052
rect 1294 3048 1298 3052
rect 1326 3048 1330 3052
rect 1454 3048 1458 3052
rect 1558 3048 1562 3052
rect 1646 3048 1650 3052
rect 1846 3048 1850 3052
rect 1918 3048 1922 3052
rect 2230 3048 2234 3052
rect 2286 3048 2290 3052
rect 2422 3048 2426 3052
rect 2430 3048 2434 3052
rect 2478 3048 2482 3052
rect 2590 3048 2594 3052
rect 3054 3048 3058 3052
rect 3358 3048 3362 3052
rect 206 3038 210 3042
rect 238 3038 242 3042
rect 718 3038 722 3042
rect 950 3038 954 3042
rect 1310 3038 1314 3042
rect 1614 3038 1618 3042
rect 1382 3028 1386 3032
rect 1862 3028 1866 3032
rect 22 3018 26 3022
rect 38 3018 42 3022
rect 46 3018 50 3022
rect 670 3018 674 3022
rect 726 3018 730 3022
rect 742 3018 746 3022
rect 766 3018 770 3022
rect 974 3018 978 3022
rect 1110 3018 1114 3022
rect 1278 3018 1282 3022
rect 1358 3018 1362 3022
rect 1430 3018 1434 3022
rect 1710 3018 1714 3022
rect 1774 3018 1778 3022
rect 1838 3018 1842 3022
rect 2254 3018 2258 3022
rect 2278 3018 2282 3022
rect 2686 3018 2690 3022
rect 2782 3018 2786 3022
rect 2798 3018 2802 3022
rect 2982 3018 2986 3022
rect 3486 3018 3490 3022
rect 3518 3018 3522 3022
rect 482 3003 486 3007
rect 489 3003 493 3007
rect 1514 3003 1518 3007
rect 1521 3003 1525 3007
rect 2538 3003 2542 3007
rect 2545 3003 2549 3007
rect 174 2988 178 2992
rect 286 2988 290 2992
rect 350 2988 354 2992
rect 462 2988 466 2992
rect 518 2988 522 2992
rect 782 2988 786 2992
rect 918 2988 922 2992
rect 966 2988 970 2992
rect 1118 2988 1122 2992
rect 1478 2988 1482 2992
rect 1582 2988 1586 2992
rect 1798 2988 1802 2992
rect 1902 2988 1906 2992
rect 2046 2988 2050 2992
rect 2102 2988 2106 2992
rect 2430 2988 2434 2992
rect 2526 2988 2530 2992
rect 2718 2988 2722 2992
rect 2750 2988 2754 2992
rect 2846 2988 2850 2992
rect 2950 2988 2954 2992
rect 2982 2988 2986 2992
rect 3126 2988 3130 2992
rect 3222 2988 3226 2992
rect 3358 2988 3362 2992
rect 1350 2978 1354 2982
rect 1446 2978 1450 2982
rect 134 2968 138 2972
rect 886 2968 890 2972
rect 1302 2968 1306 2972
rect 1862 2968 1866 2972
rect 1990 2968 1994 2972
rect 2558 2968 2562 2972
rect 3470 2968 3474 2972
rect 270 2958 274 2962
rect 366 2958 370 2962
rect 670 2958 674 2962
rect 686 2958 690 2962
rect 766 2958 770 2962
rect 790 2958 794 2962
rect 838 2958 842 2962
rect 1102 2958 1106 2962
rect 1134 2958 1138 2962
rect 1254 2958 1258 2962
rect 1286 2958 1290 2962
rect 1318 2958 1322 2962
rect 1334 2958 1338 2962
rect 1438 2958 1442 2962
rect 1526 2958 1530 2962
rect 1598 2958 1602 2962
rect 1894 2958 1898 2962
rect 1926 2958 1930 2962
rect 1982 2958 1986 2962
rect 2038 2958 2042 2962
rect 2062 2958 2066 2962
rect 2118 2958 2122 2962
rect 2158 2958 2162 2962
rect 2174 2958 2178 2962
rect 2190 2958 2194 2962
rect 2222 2958 2226 2962
rect 2302 2958 2306 2962
rect 2326 2958 2330 2962
rect 2462 2958 2466 2962
rect 2542 2958 2546 2962
rect 2830 2958 2834 2962
rect 2870 2958 2874 2962
rect 2934 2958 2938 2962
rect 2966 2958 2970 2962
rect 54 2948 58 2952
rect 78 2948 82 2952
rect 86 2948 90 2952
rect 134 2948 138 2952
rect 158 2948 162 2952
rect 38 2938 42 2942
rect 94 2938 98 2942
rect 190 2948 194 2952
rect 230 2948 234 2952
rect 262 2948 266 2952
rect 310 2948 314 2952
rect 350 2948 354 2952
rect 374 2948 378 2952
rect 390 2948 394 2952
rect 406 2948 410 2952
rect 438 2948 442 2952
rect 446 2948 450 2952
rect 470 2948 474 2952
rect 542 2948 546 2952
rect 558 2948 562 2952
rect 182 2938 186 2942
rect 254 2938 258 2942
rect 294 2938 298 2942
rect 342 2938 346 2942
rect 382 2938 386 2942
rect 638 2948 642 2952
rect 702 2948 706 2952
rect 726 2948 730 2952
rect 742 2948 746 2952
rect 846 2948 850 2952
rect 878 2948 882 2952
rect 918 2948 922 2952
rect 942 2948 946 2952
rect 990 2948 994 2952
rect 1014 2948 1018 2952
rect 1046 2948 1050 2952
rect 1062 2948 1066 2952
rect 1078 2948 1082 2952
rect 1094 2948 1098 2952
rect 1118 2948 1122 2952
rect 1158 2948 1162 2952
rect 1190 2948 1194 2952
rect 1222 2948 1226 2952
rect 1246 2948 1250 2952
rect 1254 2948 1258 2952
rect 1310 2948 1314 2952
rect 1350 2948 1354 2952
rect 1422 2948 1426 2952
rect 1558 2948 1562 2952
rect 1614 2948 1618 2952
rect 1702 2948 1706 2952
rect 1726 2948 1730 2952
rect 1742 2948 1746 2952
rect 1766 2948 1770 2952
rect 1774 2948 1778 2952
rect 1830 2948 1834 2952
rect 1838 2948 1842 2952
rect 1878 2948 1882 2952
rect 1894 2948 1898 2952
rect 1918 2948 1922 2952
rect 1950 2948 1954 2952
rect 2014 2948 2018 2952
rect 2054 2948 2058 2952
rect 2078 2948 2082 2952
rect 2102 2948 2106 2952
rect 2126 2948 2130 2952
rect 2142 2948 2146 2952
rect 2174 2948 2178 2952
rect 2206 2948 2210 2952
rect 2270 2948 2274 2952
rect 502 2938 506 2942
rect 590 2938 594 2942
rect 606 2938 610 2942
rect 622 2938 626 2942
rect 630 2938 634 2942
rect 694 2938 698 2942
rect 710 2938 714 2942
rect 734 2938 738 2942
rect 750 2938 754 2942
rect 814 2938 818 2942
rect 822 2938 826 2942
rect 838 2938 842 2942
rect 870 2938 874 2942
rect 950 2938 954 2942
rect 1022 2938 1026 2942
rect 1038 2938 1042 2942
rect 1070 2938 1074 2942
rect 1126 2938 1130 2942
rect 1150 2938 1154 2942
rect 1166 2938 1170 2942
rect 1198 2938 1202 2942
rect 1214 2938 1218 2942
rect 1278 2938 1282 2942
rect 1302 2938 1306 2942
rect 1358 2938 1362 2942
rect 1398 2938 1402 2942
rect 1430 2938 1434 2942
rect 1454 2938 1458 2942
rect 1534 2938 1538 2942
rect 1550 2938 1554 2942
rect 1566 2938 1570 2942
rect 1622 2938 1626 2942
rect 1630 2938 1634 2942
rect 1734 2938 1738 2942
rect 1766 2938 1770 2942
rect 1782 2938 1786 2942
rect 1822 2938 1826 2942
rect 1846 2938 1850 2942
rect 1870 2938 1874 2942
rect 2366 2947 2370 2951
rect 2454 2948 2458 2952
rect 2478 2948 2482 2952
rect 2518 2948 2522 2952
rect 2526 2948 2530 2952
rect 2606 2948 2610 2952
rect 2686 2948 2690 2952
rect 2710 2948 2714 2952
rect 2734 2948 2738 2952
rect 2846 2948 2850 2952
rect 2878 2948 2882 2952
rect 2902 2948 2906 2952
rect 2910 2948 2914 2952
rect 2950 2948 2954 2952
rect 2982 2948 2986 2952
rect 3006 2958 3010 2962
rect 3046 2958 3050 2962
rect 3086 2958 3090 2962
rect 3182 2958 3186 2962
rect 3238 2958 3242 2962
rect 3118 2948 3122 2952
rect 3150 2948 3154 2952
rect 3174 2948 3178 2952
rect 3190 2948 3194 2952
rect 3198 2948 3202 2952
rect 3222 2948 3226 2952
rect 3246 2948 3250 2952
rect 3262 2948 3266 2952
rect 3278 2948 3282 2952
rect 3310 2948 3314 2952
rect 1926 2938 1930 2942
rect 1958 2938 1962 2942
rect 1982 2938 1986 2942
rect 2006 2938 2010 2942
rect 2038 2938 2042 2942
rect 2054 2938 2058 2942
rect 2086 2938 2090 2942
rect 2094 2938 2098 2942
rect 2134 2938 2138 2942
rect 2182 2938 2186 2942
rect 2214 2938 2218 2942
rect 2238 2938 2242 2942
rect 2318 2938 2322 2942
rect 2374 2938 2378 2942
rect 2438 2938 2442 2942
rect 2486 2938 2490 2942
rect 2518 2938 2522 2942
rect 2646 2938 2650 2942
rect 2806 2938 2810 2942
rect 2814 2938 2818 2942
rect 2854 2938 2858 2942
rect 2918 2938 2922 2942
rect 2942 2938 2946 2942
rect 2974 2938 2978 2942
rect 3022 2938 3026 2942
rect 3030 2938 3034 2942
rect 3070 2938 3074 2942
rect 3086 2938 3090 2942
rect 3126 2938 3130 2942
rect 3142 2938 3146 2942
rect 3158 2938 3162 2942
rect 3206 2938 3210 2942
rect 3214 2938 3218 2942
rect 3254 2938 3258 2942
rect 3334 2948 3338 2952
rect 3430 2948 3434 2952
rect 3478 2948 3482 2952
rect 3518 2948 3522 2952
rect 3550 2948 3554 2952
rect 3422 2938 3426 2942
rect 6 2928 10 2932
rect 38 2928 42 2932
rect 62 2928 66 2932
rect 110 2928 114 2932
rect 118 2928 122 2932
rect 142 2928 146 2932
rect 166 2928 170 2932
rect 190 2928 194 2932
rect 206 2928 210 2932
rect 214 2928 218 2932
rect 334 2928 338 2932
rect 398 2928 402 2932
rect 406 2928 410 2932
rect 430 2928 434 2932
rect 454 2928 458 2932
rect 478 2928 482 2932
rect 566 2928 570 2932
rect 582 2928 586 2932
rect 606 2928 610 2932
rect 678 2928 682 2932
rect 718 2928 722 2932
rect 774 2928 778 2932
rect 790 2928 794 2932
rect 838 2928 842 2932
rect 886 2928 890 2932
rect 902 2928 906 2932
rect 918 2928 922 2932
rect 926 2928 930 2932
rect 966 2928 970 2932
rect 974 2928 978 2932
rect 1054 2928 1058 2932
rect 1078 2928 1082 2932
rect 1174 2928 1178 2932
rect 1182 2928 1186 2932
rect 1206 2928 1210 2932
rect 1230 2928 1234 2932
rect 1326 2928 1330 2932
rect 1374 2928 1378 2932
rect 1462 2928 1466 2932
rect 1494 2928 1498 2932
rect 1686 2928 1690 2932
rect 1798 2928 1802 2932
rect 1806 2928 1810 2932
rect 1862 2928 1866 2932
rect 1990 2928 1994 2932
rect 2150 2928 2154 2932
rect 2246 2928 2250 2932
rect 2278 2928 2282 2932
rect 2326 2928 2330 2932
rect 2454 2928 2458 2932
rect 2494 2928 2498 2932
rect 2662 2928 2666 2932
rect 2686 2928 2690 2932
rect 2862 2928 2866 2932
rect 2886 2928 2890 2932
rect 2934 2928 2938 2932
rect 3054 2928 3058 2932
rect 3094 2928 3098 2932
rect 3102 2928 3106 2932
rect 3126 2928 3130 2932
rect 3158 2928 3162 2932
rect 3270 2928 3274 2932
rect 3294 2928 3298 2932
rect 3310 2928 3314 2932
rect 3350 2928 3354 2932
rect 3374 2928 3378 2932
rect 3478 2928 3482 2932
rect 3502 2928 3506 2932
rect 3518 2928 3522 2932
rect 14 2918 18 2922
rect 70 2918 74 2922
rect 102 2918 106 2922
rect 150 2918 154 2922
rect 246 2918 250 2922
rect 326 2918 330 2922
rect 574 2918 578 2922
rect 598 2918 602 2922
rect 654 2918 658 2922
rect 766 2918 770 2922
rect 854 2918 858 2922
rect 894 2918 898 2922
rect 982 2918 986 2922
rect 1030 2918 1034 2922
rect 1238 2918 1242 2922
rect 1366 2918 1370 2922
rect 1406 2918 1410 2922
rect 1502 2918 1506 2922
rect 1598 2918 1602 2922
rect 1662 2918 1666 2922
rect 1694 2918 1698 2922
rect 1718 2918 1722 2922
rect 1742 2918 1746 2922
rect 1814 2918 1818 2922
rect 1934 2918 1938 2922
rect 2062 2918 2066 2922
rect 2190 2918 2194 2922
rect 2230 2918 2234 2922
rect 2254 2918 2258 2922
rect 2286 2918 2290 2922
rect 2310 2918 2314 2922
rect 2502 2918 2506 2922
rect 2670 2918 2674 2922
rect 2694 2918 2698 2922
rect 2718 2918 2722 2922
rect 2750 2918 2754 2922
rect 2822 2918 2826 2922
rect 3510 2918 3514 2922
rect 3534 2918 3538 2922
rect 994 2903 998 2907
rect 1001 2903 1005 2907
rect 2026 2903 2030 2907
rect 2033 2903 2037 2907
rect 3042 2903 3046 2907
rect 3049 2903 3053 2907
rect 14 2888 18 2892
rect 54 2888 58 2892
rect 78 2888 82 2892
rect 278 2888 282 2892
rect 350 2888 354 2892
rect 566 2888 570 2892
rect 590 2888 594 2892
rect 686 2888 690 2892
rect 750 2888 754 2892
rect 798 2888 802 2892
rect 1022 2888 1026 2892
rect 1046 2888 1050 2892
rect 1158 2888 1162 2892
rect 1198 2888 1202 2892
rect 1222 2888 1226 2892
rect 1294 2888 1298 2892
rect 1334 2888 1338 2892
rect 1358 2888 1362 2892
rect 1414 2888 1418 2892
rect 1558 2888 1562 2892
rect 1838 2888 1842 2892
rect 1870 2888 1874 2892
rect 1894 2888 1898 2892
rect 1918 2888 1922 2892
rect 2246 2888 2250 2892
rect 2374 2888 2378 2892
rect 2486 2888 2490 2892
rect 2518 2888 2522 2892
rect 2622 2888 2626 2892
rect 2758 2888 2762 2892
rect 2774 2888 2778 2892
rect 2870 2888 2874 2892
rect 2886 2888 2890 2892
rect 3078 2888 3082 2892
rect 3254 2888 3258 2892
rect 3398 2888 3402 2892
rect 3430 2888 3434 2892
rect 3534 2888 3538 2892
rect 6 2878 10 2882
rect 22 2878 26 2882
rect 70 2878 74 2882
rect 86 2878 90 2882
rect 94 2878 98 2882
rect 110 2878 114 2882
rect 190 2878 194 2882
rect 198 2878 202 2882
rect 230 2878 234 2882
rect 238 2878 242 2882
rect 286 2878 290 2882
rect 294 2878 298 2882
rect 302 2878 306 2882
rect 430 2878 434 2882
rect 446 2878 450 2882
rect 470 2878 474 2882
rect 558 2878 562 2882
rect 654 2878 658 2882
rect 694 2878 698 2882
rect 710 2878 714 2882
rect 742 2878 746 2882
rect 774 2878 778 2882
rect 790 2878 794 2882
rect 814 2878 818 2882
rect 830 2878 834 2882
rect 982 2878 986 2882
rect 1038 2878 1042 2882
rect 1070 2878 1074 2882
rect 1102 2878 1106 2882
rect 1150 2878 1154 2882
rect 1254 2878 1258 2882
rect 1270 2878 1274 2882
rect 1278 2878 1282 2882
rect 1350 2878 1354 2882
rect 1406 2878 1410 2882
rect 1454 2878 1458 2882
rect 1486 2878 1490 2882
rect 1550 2878 1554 2882
rect 1686 2878 1690 2882
rect 1710 2878 1714 2882
rect 1742 2878 1746 2882
rect 1846 2878 1850 2882
rect 1878 2878 1882 2882
rect 1886 2878 1890 2882
rect 1910 2878 1914 2882
rect 1950 2878 1954 2882
rect 2150 2878 2154 2882
rect 2198 2878 2202 2882
rect 2286 2878 2290 2882
rect 2390 2878 2394 2882
rect 2398 2878 2402 2882
rect 2446 2878 2450 2882
rect 2526 2878 2530 2882
rect 2598 2878 2602 2882
rect 2630 2878 2634 2882
rect 2766 2878 2770 2882
rect 2926 2878 2930 2882
rect 2958 2878 2962 2882
rect 3030 2878 3034 2882
rect 3102 2878 3106 2882
rect 3190 2878 3194 2882
rect 3238 2878 3242 2882
rect 3262 2878 3266 2882
rect 3318 2878 3322 2882
rect 3350 2878 3354 2882
rect 3382 2878 3386 2882
rect 142 2868 146 2872
rect 158 2868 162 2872
rect 230 2868 234 2872
rect 318 2868 322 2872
rect 326 2868 330 2872
rect 382 2868 386 2872
rect 422 2868 426 2872
rect 70 2858 74 2862
rect 110 2858 114 2862
rect 134 2858 138 2862
rect 166 2858 170 2862
rect 174 2858 178 2862
rect 214 2858 218 2862
rect 254 2858 258 2862
rect 262 2858 266 2862
rect 334 2858 338 2862
rect 374 2858 378 2862
rect 398 2858 402 2862
rect 414 2858 418 2862
rect 446 2858 450 2862
rect 454 2858 458 2862
rect 478 2858 482 2862
rect 510 2858 514 2862
rect 550 2868 554 2872
rect 574 2868 578 2872
rect 614 2868 618 2872
rect 646 2868 650 2872
rect 670 2868 674 2872
rect 718 2868 722 2872
rect 734 2868 738 2872
rect 806 2868 810 2872
rect 862 2868 866 2872
rect 870 2868 874 2872
rect 902 2868 906 2872
rect 934 2868 938 2872
rect 966 2868 970 2872
rect 1014 2868 1018 2872
rect 1030 2868 1034 2872
rect 1054 2868 1058 2872
rect 1102 2868 1106 2872
rect 1110 2868 1114 2872
rect 1142 2868 1146 2872
rect 1174 2868 1178 2872
rect 1206 2868 1210 2872
rect 1230 2868 1234 2872
rect 1246 2868 1250 2872
rect 1318 2868 1322 2872
rect 1326 2868 1330 2872
rect 1374 2868 1378 2872
rect 1406 2868 1410 2872
rect 1422 2868 1426 2872
rect 1430 2868 1434 2872
rect 1470 2868 1474 2872
rect 1486 2868 1490 2872
rect 1494 2868 1498 2872
rect 1566 2868 1570 2872
rect 1630 2868 1634 2872
rect 1646 2868 1650 2872
rect 1702 2868 1706 2872
rect 1726 2868 1730 2872
rect 1766 2868 1770 2872
rect 1782 2868 1786 2872
rect 1814 2868 1818 2872
rect 1830 2868 1834 2872
rect 1846 2868 1850 2872
rect 1926 2868 1930 2872
rect 1966 2868 1970 2872
rect 1974 2868 1978 2872
rect 2006 2868 2010 2872
rect 2038 2868 2042 2872
rect 2054 2868 2058 2872
rect 2094 2868 2098 2872
rect 2102 2868 2106 2872
rect 2118 2868 2122 2872
rect 2158 2868 2162 2872
rect 2206 2868 2210 2872
rect 2222 2868 2226 2872
rect 2238 2868 2242 2872
rect 2254 2868 2258 2872
rect 542 2858 546 2862
rect 582 2858 586 2862
rect 638 2858 642 2862
rect 710 2858 714 2862
rect 766 2858 770 2862
rect 774 2858 778 2862
rect 814 2858 818 2862
rect 854 2858 858 2862
rect 878 2858 882 2862
rect 894 2858 898 2862
rect 926 2858 930 2862
rect 934 2858 938 2862
rect 998 2858 1002 2862
rect 1070 2858 1074 2862
rect 1086 2858 1090 2862
rect 1118 2858 1122 2862
rect 1134 2858 1138 2862
rect 1174 2858 1178 2862
rect 1198 2858 1202 2862
rect 1230 2858 1234 2862
rect 1270 2858 1274 2862
rect 1310 2858 1314 2862
rect 1366 2858 1370 2862
rect 1382 2858 1386 2862
rect 1430 2858 1434 2862
rect 1462 2858 1466 2862
rect 1494 2858 1498 2862
rect 1526 2858 1530 2862
rect 1574 2858 1578 2862
rect 1638 2858 1642 2862
rect 1670 2858 1674 2862
rect 1718 2858 1722 2862
rect 1734 2858 1738 2862
rect 1774 2858 1778 2862
rect 1806 2858 1810 2862
rect 1822 2858 1826 2862
rect 1854 2858 1858 2862
rect 1902 2858 1906 2862
rect 1966 2858 1970 2862
rect 1982 2858 1986 2862
rect 1998 2858 2002 2862
rect 2014 2858 2018 2862
rect 2070 2858 2074 2862
rect 2118 2858 2122 2862
rect 2214 2858 2218 2862
rect 2278 2858 2282 2862
rect 2286 2858 2290 2862
rect 2302 2858 2306 2862
rect 2326 2858 2330 2862
rect 2382 2868 2386 2872
rect 2406 2868 2410 2872
rect 2430 2868 2434 2872
rect 2454 2868 2458 2872
rect 2478 2868 2482 2872
rect 2494 2868 2498 2872
rect 2502 2868 2506 2872
rect 2534 2868 2538 2872
rect 2566 2868 2570 2872
rect 2614 2868 2618 2872
rect 2638 2868 2642 2872
rect 2646 2868 2650 2872
rect 2702 2868 2706 2872
rect 2726 2868 2730 2872
rect 2734 2868 2738 2872
rect 2790 2868 2794 2872
rect 2838 2868 2842 2872
rect 2846 2868 2850 2872
rect 2854 2866 2858 2870
rect 2878 2868 2882 2872
rect 2998 2868 3002 2872
rect 3014 2868 3018 2872
rect 3054 2868 3058 2872
rect 3118 2868 3122 2872
rect 3126 2868 3130 2872
rect 3182 2868 3186 2872
rect 3206 2868 3210 2872
rect 3222 2868 3226 2872
rect 3270 2868 3274 2872
rect 3286 2868 3290 2872
rect 3318 2868 3322 2872
rect 3358 2868 3362 2872
rect 3438 2878 3442 2882
rect 3446 2878 3450 2882
rect 3486 2878 3490 2882
rect 3526 2878 3530 2882
rect 3422 2868 3426 2872
rect 3470 2868 3474 2872
rect 3494 2868 3498 2872
rect 3526 2868 3530 2872
rect 3542 2868 3546 2872
rect 2358 2858 2362 2862
rect 2414 2858 2418 2862
rect 2422 2858 2426 2862
rect 2462 2858 2466 2862
rect 2502 2858 2506 2862
rect 2558 2858 2562 2862
rect 2582 2858 2586 2862
rect 2606 2858 2610 2862
rect 2686 2858 2690 2862
rect 2718 2858 2722 2862
rect 2742 2858 2746 2862
rect 2782 2858 2786 2862
rect 2806 2858 2810 2862
rect 2830 2858 2834 2862
rect 2934 2858 2938 2862
rect 3062 2858 3066 2862
rect 3086 2858 3090 2862
rect 3190 2858 3194 2862
rect 3206 2858 3210 2862
rect 3214 2858 3218 2862
rect 3246 2858 3250 2862
rect 3262 2858 3266 2862
rect 3294 2858 3298 2862
rect 3334 2858 3338 2862
rect 3358 2858 3362 2862
rect 3406 2858 3410 2862
rect 3414 2858 3418 2862
rect 3470 2858 3474 2862
rect 3502 2858 3506 2862
rect 3550 2858 3554 2862
rect 118 2848 122 2852
rect 150 2848 154 2852
rect 198 2848 202 2852
rect 278 2848 282 2852
rect 350 2848 354 2852
rect 358 2848 362 2852
rect 414 2848 418 2852
rect 494 2848 498 2852
rect 590 2848 594 2852
rect 622 2848 626 2852
rect 670 2848 674 2852
rect 686 2848 690 2852
rect 718 2848 722 2852
rect 838 2848 842 2852
rect 910 2848 914 2852
rect 942 2848 946 2852
rect 1078 2848 1082 2852
rect 1214 2848 1218 2852
rect 1342 2848 1346 2852
rect 1398 2848 1402 2852
rect 1614 2848 1618 2852
rect 1662 2848 1666 2852
rect 1758 2848 1762 2852
rect 1790 2848 1794 2852
rect 1926 2848 1930 2852
rect 1942 2848 1946 2852
rect 2070 2848 2074 2852
rect 2174 2848 2178 2852
rect 2230 2848 2234 2852
rect 2278 2848 2282 2852
rect 2334 2848 2338 2852
rect 2366 2848 2370 2852
rect 2446 2848 2450 2852
rect 2478 2848 2482 2852
rect 2574 2848 2578 2852
rect 2694 2848 2698 2852
rect 2702 2848 2706 2852
rect 2814 2848 2818 2852
rect 3014 2848 3018 2852
rect 3110 2848 3114 2852
rect 3150 2848 3154 2852
rect 3350 2848 3354 2852
rect 3446 2848 3450 2852
rect 3518 2848 3522 2852
rect 302 2838 306 2842
rect 1294 2838 1298 2842
rect 1438 2838 1442 2842
rect 1742 2838 1746 2842
rect 2054 2838 2058 2842
rect 2318 2838 2322 2842
rect 2662 2838 2666 2842
rect 2678 2838 2682 2842
rect 2806 2838 2810 2842
rect 3054 2838 3058 2842
rect 3318 2838 3322 2842
rect 926 2828 930 2832
rect 2166 2828 2170 2832
rect 2686 2828 2690 2832
rect 134 2818 138 2822
rect 374 2818 378 2822
rect 510 2818 514 2822
rect 638 2818 642 2822
rect 798 2818 802 2822
rect 854 2818 858 2822
rect 894 2818 898 2822
rect 1134 2818 1138 2822
rect 1270 2818 1274 2822
rect 1542 2818 1546 2822
rect 1694 2818 1698 2822
rect 1806 2818 1810 2822
rect 1998 2818 2002 2822
rect 2086 2818 2090 2822
rect 2190 2818 2194 2822
rect 2326 2818 2330 2822
rect 2590 2818 2594 2822
rect 2830 2818 2834 2822
rect 2990 2818 2994 2822
rect 3094 2818 3098 2822
rect 3174 2818 3178 2822
rect 3238 2818 3242 2822
rect 3478 2818 3482 2822
rect 482 2803 486 2807
rect 489 2803 493 2807
rect 1514 2803 1518 2807
rect 1521 2803 1525 2807
rect 2538 2803 2542 2807
rect 2545 2803 2549 2807
rect 14 2788 18 2792
rect 30 2788 34 2792
rect 94 2788 98 2792
rect 118 2788 122 2792
rect 326 2788 330 2792
rect 406 2788 410 2792
rect 590 2788 594 2792
rect 614 2788 618 2792
rect 654 2788 658 2792
rect 998 2788 1002 2792
rect 1094 2788 1098 2792
rect 1134 2788 1138 2792
rect 1198 2788 1202 2792
rect 1294 2788 1298 2792
rect 1390 2788 1394 2792
rect 1486 2788 1490 2792
rect 2022 2788 2026 2792
rect 2302 2788 2306 2792
rect 2366 2788 2370 2792
rect 2438 2788 2442 2792
rect 2486 2788 2490 2792
rect 2566 2788 2570 2792
rect 2790 2788 2794 2792
rect 3030 2788 3034 2792
rect 3318 2788 3322 2792
rect 3334 2788 3338 2792
rect 3502 2788 3506 2792
rect 1574 2778 1578 2782
rect 950 2768 954 2772
rect 990 2768 994 2772
rect 1086 2768 1090 2772
rect 2110 2768 2114 2772
rect 3022 2768 3026 2772
rect 3470 2768 3474 2772
rect 3534 2768 3538 2772
rect 46 2758 50 2762
rect 78 2758 82 2762
rect 158 2758 162 2762
rect 198 2758 202 2762
rect 270 2758 274 2762
rect 774 2758 778 2762
rect 838 2758 842 2762
rect 950 2758 954 2762
rect 1006 2758 1010 2762
rect 1102 2758 1106 2762
rect 1126 2758 1130 2762
rect 1326 2758 1330 2762
rect 1430 2758 1434 2762
rect 1534 2758 1538 2762
rect 1606 2758 1610 2762
rect 30 2748 34 2752
rect 62 2748 66 2752
rect 142 2748 146 2752
rect 158 2748 162 2752
rect 198 2748 202 2752
rect 246 2748 250 2752
rect 270 2748 274 2752
rect 278 2748 282 2752
rect 302 2748 306 2752
rect 334 2748 338 2752
rect 350 2748 354 2752
rect 382 2748 386 2752
rect 454 2748 458 2752
rect 494 2748 498 2752
rect 550 2748 554 2752
rect 566 2748 570 2752
rect 670 2748 674 2752
rect 718 2748 722 2752
rect 758 2748 762 2752
rect 766 2748 770 2752
rect 782 2748 786 2752
rect 814 2748 818 2752
rect 822 2748 826 2752
rect 854 2748 858 2752
rect 870 2748 874 2752
rect 910 2748 914 2752
rect 942 2748 946 2752
rect 958 2748 962 2752
rect 998 2748 1002 2752
rect 1070 2748 1074 2752
rect 1094 2748 1098 2752
rect 1150 2748 1154 2752
rect 1182 2748 1186 2752
rect 1198 2748 1202 2752
rect 1230 2747 1234 2751
rect 1350 2748 1354 2752
rect 1382 2748 1386 2752
rect 1406 2748 1410 2752
rect 1446 2748 1450 2752
rect 1470 2748 1474 2752
rect 1566 2748 1570 2752
rect 1694 2758 1698 2762
rect 1806 2758 1810 2762
rect 1822 2758 1826 2762
rect 1886 2758 1890 2762
rect 1966 2758 1970 2762
rect 2166 2758 2170 2762
rect 2182 2758 2186 2762
rect 2214 2758 2218 2762
rect 2222 2758 2226 2762
rect 2286 2758 2290 2762
rect 2470 2758 2474 2762
rect 2502 2758 2506 2762
rect 2550 2758 2554 2762
rect 2686 2758 2690 2762
rect 1630 2748 1634 2752
rect 1710 2748 1714 2752
rect 1782 2748 1786 2752
rect 1798 2748 1802 2752
rect 1854 2748 1858 2752
rect 1870 2748 1874 2752
rect 1910 2748 1914 2752
rect 1926 2748 1930 2752
rect 1966 2748 1970 2752
rect 1974 2748 1978 2752
rect 2054 2748 2058 2752
rect 2062 2748 2066 2752
rect 2110 2748 2114 2752
rect 2190 2748 2194 2752
rect 2222 2748 2226 2752
rect 2238 2748 2242 2752
rect 2262 2748 2266 2752
rect 2278 2748 2282 2752
rect 2302 2748 2306 2752
rect 2358 2748 2362 2752
rect 2414 2748 2418 2752
rect 2462 2748 2466 2752
rect 2486 2748 2490 2752
rect 2518 2748 2522 2752
rect 2550 2748 2554 2752
rect 2566 2748 2570 2752
rect 2582 2748 2586 2752
rect 2630 2748 2634 2752
rect 2638 2748 2642 2752
rect 2654 2748 2658 2752
rect 2670 2748 2674 2752
rect 2750 2748 2754 2752
rect 2798 2748 2802 2752
rect 2814 2748 2818 2752
rect 2926 2758 2930 2762
rect 2998 2758 3002 2762
rect 3038 2758 3042 2762
rect 3142 2758 3146 2762
rect 3198 2758 3202 2762
rect 3262 2758 3266 2762
rect 3286 2758 3290 2762
rect 3398 2758 3402 2762
rect 3430 2758 3434 2762
rect 2894 2748 2898 2752
rect 2966 2748 2970 2752
rect 2974 2748 2978 2752
rect 3006 2748 3010 2752
rect 3030 2748 3034 2752
rect 3070 2748 3074 2752
rect 3086 2748 3090 2752
rect 3134 2748 3138 2752
rect 3158 2748 3162 2752
rect 3182 2748 3186 2752
rect 3230 2748 3234 2752
rect 3254 2748 3258 2752
rect 3278 2748 3282 2752
rect 3302 2748 3306 2752
rect 3382 2748 3386 2752
rect 3406 2748 3410 2752
rect 3414 2748 3418 2752
rect 3422 2748 3426 2752
rect 3446 2748 3450 2752
rect 3486 2748 3490 2752
rect 3502 2748 3506 2752
rect 3542 2748 3546 2752
rect 6 2738 10 2742
rect 22 2738 26 2742
rect 54 2738 58 2742
rect 134 2738 138 2742
rect 158 2738 162 2742
rect 182 2738 186 2742
rect 278 2738 282 2742
rect 294 2738 298 2742
rect 310 2738 314 2742
rect 326 2738 330 2742
rect 358 2738 362 2742
rect 414 2738 418 2742
rect 438 2738 442 2742
rect 510 2738 514 2742
rect 558 2738 562 2742
rect 582 2738 586 2742
rect 598 2738 602 2742
rect 606 2738 610 2742
rect 638 2738 642 2742
rect 678 2738 682 2742
rect 726 2738 730 2742
rect 790 2738 794 2742
rect 806 2738 810 2742
rect 846 2738 850 2742
rect 862 2738 866 2742
rect 886 2738 890 2742
rect 910 2738 914 2742
rect 934 2738 938 2742
rect 974 2738 978 2742
rect 1062 2738 1066 2742
rect 1110 2738 1114 2742
rect 1142 2738 1146 2742
rect 1158 2738 1162 2742
rect 1214 2738 1218 2742
rect 1342 2738 1346 2742
rect 1358 2738 1362 2742
rect 1374 2738 1378 2742
rect 1398 2738 1402 2742
rect 1454 2738 1458 2742
rect 1462 2738 1466 2742
rect 1582 2738 1586 2742
rect 1590 2738 1594 2742
rect 1638 2738 1642 2742
rect 1702 2738 1706 2742
rect 1774 2738 1778 2742
rect 1806 2738 1810 2742
rect 1862 2738 1866 2742
rect 1894 2738 1898 2742
rect 1918 2738 1922 2742
rect 1974 2738 1978 2742
rect 1990 2738 1994 2742
rect 2070 2738 2074 2742
rect 2118 2738 2122 2742
rect 2142 2738 2146 2742
rect 2198 2738 2202 2742
rect 2246 2738 2250 2742
rect 2270 2738 2274 2742
rect 2342 2738 2346 2742
rect 2350 2738 2354 2742
rect 2374 2738 2378 2742
rect 2382 2738 2386 2742
rect 2430 2738 2434 2742
rect 2454 2738 2458 2742
rect 2494 2738 2498 2742
rect 2526 2738 2530 2742
rect 2574 2738 2578 2742
rect 2662 2738 2666 2742
rect 2742 2738 2746 2742
rect 2758 2738 2762 2742
rect 2806 2738 2810 2742
rect 2838 2738 2842 2742
rect 2854 2738 2858 2742
rect 2918 2738 2922 2742
rect 2942 2738 2946 2742
rect 2982 2738 2986 2742
rect 2998 2738 3002 2742
rect 3078 2738 3082 2742
rect 3110 2738 3114 2742
rect 3166 2738 3170 2742
rect 3174 2738 3178 2742
rect 3190 2738 3194 2742
rect 3222 2738 3226 2742
rect 3278 2738 3282 2742
rect 3310 2738 3314 2742
rect 3350 2740 3354 2744
rect 3358 2738 3362 2742
rect 3390 2738 3394 2742
rect 3422 2738 3426 2742
rect 3454 2738 3458 2742
rect 3510 2738 3514 2742
rect 3518 2740 3522 2744
rect 3558 2738 3562 2742
rect 206 2728 210 2732
rect 222 2728 226 2732
rect 230 2728 234 2732
rect 326 2728 330 2732
rect 350 2728 354 2732
rect 398 2728 402 2732
rect 422 2728 426 2732
rect 478 2728 482 2732
rect 526 2728 530 2732
rect 534 2728 538 2732
rect 582 2728 586 2732
rect 622 2728 626 2732
rect 662 2728 666 2732
rect 694 2728 698 2732
rect 702 2728 706 2732
rect 710 2728 714 2732
rect 742 2728 746 2732
rect 806 2728 810 2732
rect 838 2728 842 2732
rect 886 2728 890 2732
rect 918 2728 922 2732
rect 1030 2728 1034 2732
rect 1174 2728 1178 2732
rect 1182 2728 1186 2732
rect 1302 2728 1306 2732
rect 1318 2728 1322 2732
rect 1334 2728 1338 2732
rect 1422 2728 1426 2732
rect 1494 2728 1498 2732
rect 1534 2728 1538 2732
rect 1550 2728 1554 2732
rect 1566 2728 1570 2732
rect 1646 2728 1650 2732
rect 1678 2728 1682 2732
rect 1726 2728 1730 2732
rect 1734 2728 1738 2732
rect 1782 2728 1786 2732
rect 2006 2728 2010 2732
rect 2038 2728 2042 2732
rect 2086 2728 2090 2732
rect 2126 2728 2130 2732
rect 2174 2728 2178 2732
rect 2254 2728 2258 2732
rect 2326 2728 2330 2732
rect 2334 2728 2338 2732
rect 2438 2728 2442 2732
rect 2598 2728 2602 2732
rect 2654 2728 2658 2732
rect 2774 2728 2778 2732
rect 2782 2728 2786 2732
rect 2798 2728 2802 2732
rect 2886 2728 2890 2732
rect 2950 2728 2954 2732
rect 3054 2728 3058 2732
rect 3094 2728 3098 2732
rect 3134 2728 3138 2732
rect 3206 2728 3210 2732
rect 3238 2728 3242 2732
rect 3326 2728 3330 2732
rect 3462 2728 3466 2732
rect 3486 2728 3490 2732
rect 14 2718 18 2722
rect 190 2718 194 2722
rect 430 2718 434 2722
rect 470 2718 474 2722
rect 630 2718 634 2722
rect 686 2718 690 2722
rect 894 2718 898 2722
rect 926 2718 930 2722
rect 1054 2718 1058 2722
rect 1118 2718 1122 2722
rect 1366 2718 1370 2722
rect 1414 2718 1418 2722
rect 1430 2718 1434 2722
rect 1502 2718 1506 2722
rect 1614 2718 1618 2722
rect 1654 2718 1658 2722
rect 1718 2718 1722 2722
rect 1750 2718 1754 2722
rect 1814 2718 1818 2722
rect 1838 2718 1842 2722
rect 2166 2718 2170 2722
rect 2222 2718 2226 2722
rect 2502 2718 2506 2722
rect 2614 2718 2618 2722
rect 2726 2718 2730 2722
rect 2766 2718 2770 2722
rect 2830 2718 2834 2722
rect 2846 2718 2850 2722
rect 2870 2718 2874 2722
rect 2926 2718 2930 2722
rect 2958 2718 2962 2722
rect 3102 2718 3106 2722
rect 3142 2718 3146 2722
rect 3214 2718 3218 2722
rect 3286 2718 3290 2722
rect 3366 2718 3370 2722
rect 994 2703 998 2707
rect 1001 2703 1005 2707
rect 2026 2703 2030 2707
rect 2033 2703 2037 2707
rect 3042 2703 3046 2707
rect 3049 2703 3053 2707
rect 198 2688 202 2692
rect 222 2688 226 2692
rect 278 2688 282 2692
rect 430 2688 434 2692
rect 518 2688 522 2692
rect 550 2688 554 2692
rect 614 2688 618 2692
rect 662 2688 666 2692
rect 838 2688 842 2692
rect 926 2688 930 2692
rect 1022 2688 1026 2692
rect 1046 2688 1050 2692
rect 1166 2688 1170 2692
rect 1230 2688 1234 2692
rect 1286 2688 1290 2692
rect 1334 2688 1338 2692
rect 1398 2688 1402 2692
rect 1806 2688 1810 2692
rect 1830 2688 1834 2692
rect 1926 2688 1930 2692
rect 1982 2688 1986 2692
rect 2046 2688 2050 2692
rect 2142 2688 2146 2692
rect 2238 2688 2242 2692
rect 2430 2688 2434 2692
rect 2446 2688 2450 2692
rect 2478 2688 2482 2692
rect 2630 2688 2634 2692
rect 2646 2688 2650 2692
rect 2670 2688 2674 2692
rect 2758 2688 2762 2692
rect 2798 2688 2802 2692
rect 2830 2688 2834 2692
rect 2950 2688 2954 2692
rect 2982 2688 2986 2692
rect 3046 2688 3050 2692
rect 3134 2688 3138 2692
rect 3166 2688 3170 2692
rect 3270 2688 3274 2692
rect 3302 2688 3306 2692
rect 3318 2688 3322 2692
rect 3358 2688 3362 2692
rect 3390 2688 3394 2692
rect 3446 2688 3450 2692
rect 6 2678 10 2682
rect 62 2678 66 2682
rect 78 2678 82 2682
rect 94 2678 98 2682
rect 102 2678 106 2682
rect 190 2678 194 2682
rect 214 2678 218 2682
rect 254 2678 258 2682
rect 286 2678 290 2682
rect 350 2678 354 2682
rect 22 2668 26 2672
rect 38 2668 42 2672
rect 62 2668 66 2672
rect 126 2668 130 2672
rect 158 2668 162 2672
rect 174 2668 178 2672
rect 270 2668 274 2672
rect 286 2668 290 2672
rect 318 2668 322 2672
rect 446 2678 450 2682
rect 510 2678 514 2682
rect 670 2678 674 2682
rect 678 2678 682 2682
rect 726 2678 730 2682
rect 758 2678 762 2682
rect 774 2678 778 2682
rect 798 2678 802 2682
rect 830 2678 834 2682
rect 982 2678 986 2682
rect 1030 2678 1034 2682
rect 1110 2678 1114 2682
rect 1174 2678 1178 2682
rect 1222 2678 1226 2682
rect 1526 2678 1530 2682
rect 1646 2678 1650 2682
rect 1686 2678 1690 2682
rect 1694 2678 1698 2682
rect 1726 2678 1730 2682
rect 1838 2678 1842 2682
rect 1918 2678 1922 2682
rect 1966 2678 1970 2682
rect 2006 2678 2010 2682
rect 2070 2678 2074 2682
rect 2110 2678 2114 2682
rect 2126 2678 2130 2682
rect 2134 2678 2138 2682
rect 2214 2678 2218 2682
rect 2246 2678 2250 2682
rect 2254 2678 2258 2682
rect 2278 2678 2282 2682
rect 2302 2678 2306 2682
rect 2358 2678 2362 2682
rect 2382 2678 2386 2682
rect 2398 2678 2402 2682
rect 2438 2678 2442 2682
rect 2494 2678 2498 2682
rect 2550 2678 2554 2682
rect 2606 2678 2610 2682
rect 2638 2678 2642 2682
rect 2654 2678 2658 2682
rect 2766 2678 2770 2682
rect 2838 2678 2842 2682
rect 2846 2678 2850 2682
rect 2862 2678 2866 2682
rect 2958 2678 2962 2682
rect 2990 2678 2994 2682
rect 3174 2678 3178 2682
rect 3198 2678 3202 2682
rect 3206 2678 3210 2682
rect 3278 2678 3282 2682
rect 3366 2678 3370 2682
rect 3382 2678 3386 2682
rect 3422 2678 3426 2682
rect 3430 2678 3434 2682
rect 3438 2678 3442 2682
rect 3478 2678 3482 2682
rect 390 2668 394 2672
rect 406 2668 410 2672
rect 422 2668 426 2672
rect 526 2668 530 2672
rect 558 2668 562 2672
rect 590 2668 594 2672
rect 606 2668 610 2672
rect 638 2668 642 2672
rect 654 2668 658 2672
rect 694 2668 698 2672
rect 734 2668 738 2672
rect 758 2668 762 2672
rect 846 2668 850 2672
rect 878 2668 882 2672
rect 894 2668 898 2672
rect 950 2668 954 2672
rect 1014 2668 1018 2672
rect 1054 2668 1058 2672
rect 1078 2668 1082 2672
rect 1094 2668 1098 2672
rect 1110 2668 1114 2672
rect 1158 2668 1162 2672
rect 1238 2668 1242 2672
rect 6 2658 10 2662
rect 30 2658 34 2662
rect 46 2658 50 2662
rect 78 2658 82 2662
rect 94 2658 98 2662
rect 118 2658 122 2662
rect 166 2658 170 2662
rect 206 2658 210 2662
rect 230 2658 234 2662
rect 238 2658 242 2662
rect 262 2658 266 2662
rect 294 2658 298 2662
rect 310 2658 314 2662
rect 326 2658 330 2662
rect 334 2658 338 2662
rect 374 2658 378 2662
rect 382 2658 386 2662
rect 414 2658 418 2662
rect 462 2658 466 2662
rect 534 2658 538 2662
rect 566 2658 570 2662
rect 582 2658 586 2662
rect 630 2658 634 2662
rect 646 2658 650 2662
rect 702 2658 706 2662
rect 774 2658 778 2662
rect 782 2658 786 2662
rect 798 2658 802 2662
rect 854 2658 858 2662
rect 902 2658 906 2662
rect 942 2658 946 2662
rect 1086 2658 1090 2662
rect 1262 2666 1266 2670
rect 1270 2668 1274 2672
rect 1318 2668 1322 2672
rect 1454 2668 1458 2672
rect 1470 2668 1474 2672
rect 1510 2668 1514 2672
rect 1542 2668 1546 2672
rect 1590 2668 1594 2672
rect 1606 2668 1610 2672
rect 1614 2668 1618 2672
rect 1638 2668 1642 2672
rect 1662 2668 1666 2672
rect 1694 2668 1698 2672
rect 1766 2668 1770 2672
rect 1782 2668 1786 2672
rect 1822 2668 1826 2672
rect 1870 2668 1874 2672
rect 1894 2668 1898 2672
rect 2062 2668 2066 2672
rect 2094 2668 2098 2672
rect 2110 2668 2114 2672
rect 2150 2668 2154 2672
rect 2158 2668 2162 2672
rect 2198 2668 2202 2672
rect 2214 2668 2218 2672
rect 2230 2668 2234 2672
rect 1126 2658 1130 2662
rect 1150 2658 1154 2662
rect 1206 2658 1210 2662
rect 1238 2658 1242 2662
rect 1302 2658 1306 2662
rect 1350 2658 1354 2662
rect 1366 2658 1370 2662
rect 1414 2658 1418 2662
rect 1422 2658 1426 2662
rect 1494 2658 1498 2662
rect 1542 2658 1546 2662
rect 1558 2658 1562 2662
rect 1582 2658 1586 2662
rect 1614 2658 1618 2662
rect 1654 2658 1658 2662
rect 1670 2658 1674 2662
rect 1678 2658 1682 2662
rect 1742 2658 1746 2662
rect 1774 2658 1778 2662
rect 1790 2658 1794 2662
rect 1814 2658 1818 2662
rect 1854 2658 1858 2662
rect 1902 2658 1906 2662
rect 1918 2658 1922 2662
rect 1942 2658 1946 2662
rect 2006 2658 2010 2662
rect 2022 2658 2026 2662
rect 2110 2658 2114 2662
rect 2158 2658 2162 2662
rect 2222 2658 2226 2662
rect 2302 2658 2306 2662
rect 2318 2658 2322 2662
rect 2342 2658 2346 2662
rect 2406 2668 2410 2672
rect 2414 2666 2418 2670
rect 2470 2668 2474 2672
rect 2462 2658 2466 2662
rect 2558 2668 2562 2672
rect 2598 2668 2602 2672
rect 2622 2668 2626 2672
rect 2662 2668 2666 2672
rect 2686 2668 2690 2672
rect 2710 2668 2714 2672
rect 2734 2668 2738 2672
rect 2750 2668 2754 2672
rect 2774 2668 2778 2672
rect 2806 2668 2810 2672
rect 2822 2668 2826 2672
rect 2878 2668 2882 2672
rect 2894 2668 2898 2672
rect 2910 2668 2914 2672
rect 2926 2668 2930 2672
rect 2942 2668 2946 2672
rect 2974 2668 2978 2672
rect 3006 2668 3010 2672
rect 3030 2668 3034 2672
rect 3118 2668 3122 2672
rect 3134 2668 3138 2672
rect 3150 2668 3154 2672
rect 3246 2668 3250 2672
rect 3262 2668 3266 2672
rect 3286 2668 3290 2672
rect 3334 2668 3338 2672
rect 3350 2668 3354 2672
rect 3406 2668 3410 2672
rect 3454 2668 3458 2672
rect 3486 2668 3490 2672
rect 3494 2668 3498 2672
rect 2494 2658 2498 2662
rect 2510 2658 2514 2662
rect 2526 2658 2530 2662
rect 2534 2658 2538 2662
rect 2574 2658 2578 2662
rect 2614 2658 2618 2662
rect 2742 2658 2746 2662
rect 2782 2658 2786 2662
rect 2798 2658 2802 2662
rect 2814 2658 2818 2662
rect 2846 2658 2850 2662
rect 2870 2658 2874 2662
rect 2910 2658 2914 2662
rect 2926 2658 2930 2662
rect 2966 2658 2970 2662
rect 2998 2658 3002 2662
rect 3030 2658 3034 2662
rect 3070 2658 3074 2662
rect 3102 2658 3106 2662
rect 3158 2658 3162 2662
rect 3182 2658 3186 2662
rect 3198 2658 3202 2662
rect 3222 2658 3226 2662
rect 3246 2658 3250 2662
rect 3342 2658 3346 2662
rect 3414 2658 3418 2662
rect 150 2648 154 2652
rect 182 2648 186 2652
rect 438 2648 442 2652
rect 550 2648 554 2652
rect 614 2648 618 2652
rect 718 2648 722 2652
rect 806 2648 810 2652
rect 870 2648 874 2652
rect 918 2648 922 2652
rect 926 2648 930 2652
rect 1038 2648 1042 2652
rect 1062 2648 1066 2652
rect 1118 2648 1122 2652
rect 1182 2648 1186 2652
rect 1358 2648 1362 2652
rect 1454 2648 1458 2652
rect 1534 2648 1538 2652
rect 1574 2648 1578 2652
rect 1590 2648 1594 2652
rect 1622 2648 1626 2652
rect 1718 2648 1722 2652
rect 1846 2648 1850 2652
rect 1878 2648 1882 2652
rect 2182 2648 2186 2652
rect 2326 2648 2330 2652
rect 2470 2648 2474 2652
rect 2678 2648 2682 2652
rect 2718 2648 2722 2652
rect 2910 2648 2914 2652
rect 3086 2648 3090 2652
rect 3230 2648 3234 2652
rect 3390 2648 3394 2652
rect 118 2638 122 2642
rect 478 2638 482 2642
rect 598 2638 602 2642
rect 702 2638 706 2642
rect 774 2638 778 2642
rect 822 2638 826 2642
rect 886 2638 890 2642
rect 1118 2638 1122 2642
rect 1134 2638 1138 2642
rect 1374 2638 1378 2642
rect 2582 2638 2586 2642
rect 3510 2638 3514 2642
rect 686 2628 690 2632
rect 902 2628 906 2632
rect 1206 2628 1210 2632
rect 134 2618 138 2622
rect 390 2618 394 2622
rect 566 2618 570 2622
rect 854 2618 858 2622
rect 1070 2618 1074 2622
rect 1126 2618 1130 2622
rect 1190 2618 1194 2622
rect 1310 2618 1314 2622
rect 1382 2618 1386 2622
rect 1494 2618 1498 2622
rect 1558 2618 1562 2622
rect 1710 2618 1714 2622
rect 1750 2618 1754 2622
rect 1886 2618 1890 2622
rect 2262 2618 2266 2622
rect 2310 2618 2314 2622
rect 2342 2618 2346 2622
rect 2894 2618 2898 2622
rect 3006 2618 3010 2622
rect 3182 2618 3186 2622
rect 3238 2618 3242 2622
rect 3374 2618 3378 2622
rect 3398 2618 3402 2622
rect 3462 2618 3466 2622
rect 482 2603 486 2607
rect 489 2603 493 2607
rect 1514 2603 1518 2607
rect 1521 2603 1525 2607
rect 2538 2603 2542 2607
rect 2545 2603 2549 2607
rect 14 2588 18 2592
rect 38 2588 42 2592
rect 102 2588 106 2592
rect 174 2588 178 2592
rect 222 2588 226 2592
rect 262 2588 266 2592
rect 398 2588 402 2592
rect 598 2588 602 2592
rect 686 2588 690 2592
rect 750 2588 754 2592
rect 798 2588 802 2592
rect 830 2588 834 2592
rect 878 2588 882 2592
rect 1238 2588 1242 2592
rect 1294 2588 1298 2592
rect 1574 2588 1578 2592
rect 1814 2588 1818 2592
rect 1838 2588 1842 2592
rect 1974 2588 1978 2592
rect 2366 2588 2370 2592
rect 2382 2588 2386 2592
rect 2430 2588 2434 2592
rect 2606 2588 2610 2592
rect 2718 2588 2722 2592
rect 2854 2588 2858 2592
rect 3238 2588 3242 2592
rect 3246 2588 3250 2592
rect 3286 2588 3290 2592
rect 3406 2588 3410 2592
rect 646 2578 650 2582
rect 2582 2578 2586 2582
rect 3550 2578 3554 2582
rect 718 2568 722 2572
rect 782 2568 786 2572
rect 822 2568 826 2572
rect 1078 2568 1082 2572
rect 1278 2568 1282 2572
rect 1398 2568 1402 2572
rect 2614 2568 2618 2572
rect 2814 2568 2818 2572
rect 2958 2568 2962 2572
rect 3054 2568 3058 2572
rect 3350 2568 3354 2572
rect 54 2558 58 2562
rect 126 2558 130 2562
rect 110 2548 114 2552
rect 134 2548 138 2552
rect 190 2548 194 2552
rect 222 2548 226 2552
rect 246 2558 250 2562
rect 318 2558 322 2562
rect 454 2558 458 2562
rect 566 2558 570 2562
rect 582 2558 586 2562
rect 622 2558 626 2562
rect 702 2558 706 2562
rect 726 2558 730 2562
rect 734 2558 738 2562
rect 838 2558 842 2562
rect 870 2558 874 2562
rect 902 2558 906 2562
rect 1166 2558 1170 2562
rect 1198 2558 1202 2562
rect 1350 2558 1354 2562
rect 1478 2558 1482 2562
rect 1486 2558 1490 2562
rect 1590 2558 1594 2562
rect 1678 2558 1682 2562
rect 1694 2558 1698 2562
rect 1758 2558 1762 2562
rect 1766 2558 1770 2562
rect 1854 2558 1858 2562
rect 1958 2558 1962 2562
rect 2006 2558 2010 2562
rect 2102 2558 2106 2562
rect 2166 2558 2170 2562
rect 2190 2558 2194 2562
rect 2414 2558 2418 2562
rect 2446 2558 2450 2562
rect 262 2548 266 2552
rect 302 2548 306 2552
rect 334 2548 338 2552
rect 358 2548 362 2552
rect 374 2548 378 2552
rect 398 2548 402 2552
rect 422 2548 426 2552
rect 446 2548 450 2552
rect 470 2548 474 2552
rect 510 2548 514 2552
rect 526 2548 530 2552
rect 534 2548 538 2552
rect 2494 2558 2498 2562
rect 2566 2558 2570 2562
rect 2598 2558 2602 2562
rect 2646 2558 2650 2562
rect 2654 2558 2658 2562
rect 2734 2558 2738 2562
rect 590 2548 594 2552
rect 614 2548 618 2552
rect 710 2548 714 2552
rect 766 2548 770 2552
rect 790 2548 794 2552
rect 830 2548 834 2552
rect 934 2548 938 2552
rect 966 2548 970 2552
rect 1014 2548 1018 2552
rect 1110 2548 1114 2552
rect 1142 2548 1146 2552
rect 1174 2548 1178 2552
rect 1214 2548 1218 2552
rect 1310 2548 1314 2552
rect 1334 2548 1338 2552
rect 1366 2548 1370 2552
rect 6 2538 10 2542
rect 30 2538 34 2542
rect 70 2538 74 2542
rect 158 2538 162 2542
rect 182 2538 186 2542
rect 214 2538 218 2542
rect 270 2538 274 2542
rect 278 2538 282 2542
rect 294 2538 298 2542
rect 326 2538 330 2542
rect 478 2538 482 2542
rect 518 2538 522 2542
rect 542 2538 546 2542
rect 566 2538 570 2542
rect 758 2538 762 2542
rect 766 2538 770 2542
rect 806 2538 810 2542
rect 846 2538 850 2542
rect 894 2538 898 2542
rect 918 2538 922 2542
rect 926 2538 930 2542
rect 958 2538 962 2542
rect 1006 2538 1010 2542
rect 1046 2538 1050 2542
rect 1054 2538 1058 2542
rect 1078 2538 1082 2542
rect 1086 2540 1090 2544
rect 1118 2538 1122 2542
rect 1134 2538 1138 2542
rect 1142 2538 1146 2542
rect 1222 2538 1226 2542
rect 1230 2538 1234 2542
rect 1246 2538 1250 2542
rect 1262 2538 1266 2542
rect 1406 2538 1410 2542
rect 1462 2548 1466 2552
rect 1542 2548 1546 2552
rect 1550 2548 1554 2552
rect 1582 2548 1586 2552
rect 1606 2548 1610 2552
rect 1646 2548 1650 2552
rect 1662 2548 1666 2552
rect 1670 2548 1674 2552
rect 1702 2548 1706 2552
rect 1734 2548 1738 2552
rect 1838 2548 1842 2552
rect 1862 2548 1866 2552
rect 1878 2548 1882 2552
rect 1894 2548 1898 2552
rect 1934 2548 1938 2552
rect 1950 2548 1954 2552
rect 2014 2548 2018 2552
rect 2038 2548 2042 2552
rect 2214 2548 2218 2552
rect 2262 2548 2266 2552
rect 2286 2548 2290 2552
rect 2350 2548 2354 2552
rect 2406 2548 2410 2552
rect 2486 2548 2490 2552
rect 2510 2548 2514 2552
rect 2518 2548 2522 2552
rect 2582 2548 2586 2552
rect 2606 2548 2610 2552
rect 2670 2548 2674 2552
rect 2886 2558 2890 2562
rect 2918 2558 2922 2562
rect 2870 2548 2874 2552
rect 2894 2548 2898 2552
rect 2934 2548 2938 2552
rect 2958 2548 2962 2552
rect 2982 2558 2986 2562
rect 3094 2558 3098 2562
rect 3118 2558 3122 2562
rect 3222 2558 3226 2562
rect 3342 2558 3346 2562
rect 3366 2558 3370 2562
rect 2998 2548 3002 2552
rect 3014 2548 3018 2552
rect 3078 2548 3082 2552
rect 3134 2548 3138 2552
rect 3150 2548 3154 2552
rect 3198 2548 3202 2552
rect 3270 2548 3274 2552
rect 3278 2548 3282 2552
rect 3318 2548 3322 2552
rect 3334 2548 3338 2552
rect 3470 2548 3474 2552
rect 3486 2548 3490 2552
rect 1438 2538 1442 2542
rect 1454 2538 1458 2542
rect 1526 2538 1530 2542
rect 1542 2538 1546 2542
rect 1558 2538 1562 2542
rect 1574 2538 1578 2542
rect 1614 2538 1618 2542
rect 1638 2538 1642 2542
rect 1654 2538 1658 2542
rect 1726 2538 1730 2542
rect 1742 2538 1746 2542
rect 1766 2538 1770 2542
rect 1782 2538 1786 2542
rect 1822 2538 1826 2542
rect 1830 2538 1834 2542
rect 1870 2538 1874 2542
rect 1942 2538 1946 2542
rect 1982 2538 1986 2542
rect 1990 2538 1994 2542
rect 2014 2538 2018 2542
rect 2038 2538 2042 2542
rect 2086 2540 2090 2544
rect 2094 2538 2098 2542
rect 2126 2538 2130 2542
rect 2150 2538 2154 2542
rect 2158 2538 2162 2542
rect 2174 2538 2178 2542
rect 2190 2538 2194 2542
rect 2238 2538 2242 2542
rect 2294 2538 2298 2542
rect 2310 2538 2314 2542
rect 2342 2538 2346 2542
rect 2358 2538 2362 2542
rect 2438 2538 2442 2542
rect 2462 2538 2466 2542
rect 2470 2538 2474 2542
rect 2486 2538 2490 2542
rect 2526 2538 2530 2542
rect 2590 2538 2594 2542
rect 2630 2538 2634 2542
rect 2646 2538 2650 2542
rect 2678 2538 2682 2542
rect 2726 2538 2730 2542
rect 2750 2538 2754 2542
rect 2822 2538 2826 2542
rect 2846 2538 2850 2542
rect 2862 2538 2866 2542
rect 2942 2538 2946 2542
rect 2950 2538 2954 2542
rect 3006 2538 3010 2542
rect 3022 2538 3026 2542
rect 3094 2538 3098 2542
rect 3110 2538 3114 2542
rect 3142 2538 3146 2542
rect 3158 2538 3162 2542
rect 3206 2538 3210 2542
rect 3262 2538 3266 2542
rect 3350 2538 3354 2542
rect 3374 2538 3378 2542
rect 3422 2538 3426 2542
rect 3438 2538 3442 2542
rect 38 2528 42 2532
rect 78 2528 82 2532
rect 94 2528 98 2532
rect 110 2528 114 2532
rect 134 2528 138 2532
rect 158 2528 162 2532
rect 374 2528 378 2532
rect 382 2528 386 2532
rect 406 2528 410 2532
rect 502 2528 506 2532
rect 558 2528 562 2532
rect 606 2528 610 2532
rect 630 2528 634 2532
rect 670 2528 674 2532
rect 694 2528 698 2532
rect 870 2528 874 2532
rect 1134 2528 1138 2532
rect 1174 2528 1178 2532
rect 1318 2528 1322 2532
rect 1414 2528 1418 2532
rect 1430 2528 1434 2532
rect 1518 2528 1522 2532
rect 1622 2528 1626 2532
rect 1686 2528 1690 2532
rect 1710 2528 1714 2532
rect 1886 2528 1890 2532
rect 1910 2528 1914 2532
rect 1926 2528 1930 2532
rect 2030 2528 2034 2532
rect 2046 2528 2050 2532
rect 2062 2528 2066 2532
rect 2182 2528 2186 2532
rect 2206 2528 2210 2532
rect 2254 2528 2258 2532
rect 2326 2528 2330 2532
rect 2374 2528 2378 2532
rect 2390 2528 2394 2532
rect 2542 2528 2546 2532
rect 2686 2528 2690 2532
rect 2758 2528 2762 2532
rect 2790 2528 2794 2532
rect 2838 2528 2842 2532
rect 3038 2528 3042 2532
rect 3166 2528 3170 2532
rect 3182 2528 3186 2532
rect 3230 2528 3234 2532
rect 3246 2528 3250 2532
rect 3310 2528 3314 2532
rect 14 2518 18 2522
rect 54 2518 58 2522
rect 150 2518 154 2522
rect 174 2518 178 2522
rect 206 2518 210 2522
rect 286 2518 290 2522
rect 318 2518 322 2522
rect 350 2518 354 2522
rect 438 2518 442 2522
rect 454 2518 458 2522
rect 574 2518 578 2522
rect 774 2518 778 2522
rect 854 2518 858 2522
rect 878 2518 882 2522
rect 886 2518 890 2522
rect 910 2518 914 2522
rect 950 2518 954 2522
rect 982 2518 986 2522
rect 1030 2518 1034 2522
rect 1038 2518 1042 2522
rect 1062 2518 1066 2522
rect 1102 2518 1106 2522
rect 1182 2518 1186 2522
rect 1238 2518 1242 2522
rect 1254 2518 1258 2522
rect 1270 2518 1274 2522
rect 1326 2518 1330 2522
rect 1446 2518 1450 2522
rect 1478 2518 1482 2522
rect 1494 2518 1498 2522
rect 1590 2518 1594 2522
rect 1630 2518 1634 2522
rect 1718 2518 1722 2522
rect 1774 2518 1778 2522
rect 2070 2518 2074 2522
rect 2102 2518 2106 2522
rect 2278 2518 2282 2522
rect 2398 2518 2402 2522
rect 2486 2518 2490 2522
rect 2646 2518 2650 2522
rect 2766 2518 2770 2522
rect 2886 2518 2890 2522
rect 2902 2518 2906 2522
rect 3030 2518 3034 2522
rect 3094 2518 3098 2522
rect 3118 2518 3122 2522
rect 3286 2518 3290 2522
rect 3366 2518 3370 2522
rect 3518 2518 3522 2522
rect 994 2503 998 2507
rect 1001 2503 1005 2507
rect 2026 2503 2030 2507
rect 2033 2503 2037 2507
rect 3042 2503 3046 2507
rect 3049 2503 3053 2507
rect 46 2488 50 2492
rect 70 2488 74 2492
rect 158 2488 162 2492
rect 198 2488 202 2492
rect 222 2488 226 2492
rect 1318 2488 1322 2492
rect 1446 2488 1450 2492
rect 1630 2488 1634 2492
rect 1734 2488 1738 2492
rect 1790 2488 1794 2492
rect 1854 2488 1858 2492
rect 1958 2488 1962 2492
rect 1998 2488 2002 2492
rect 2158 2488 2162 2492
rect 2174 2488 2178 2492
rect 2206 2488 2210 2492
rect 2286 2488 2290 2492
rect 2302 2488 2306 2492
rect 2398 2488 2402 2492
rect 2414 2488 2418 2492
rect 2470 2488 2474 2492
rect 2582 2488 2586 2492
rect 2598 2488 2602 2492
rect 2806 2488 2810 2492
rect 2846 2488 2850 2492
rect 2918 2488 2922 2492
rect 3142 2488 3146 2492
rect 3158 2488 3162 2492
rect 3190 2488 3194 2492
rect 3286 2488 3290 2492
rect 3342 2488 3346 2492
rect 3470 2488 3474 2492
rect 142 2478 146 2482
rect 206 2478 210 2482
rect 230 2478 234 2482
rect 342 2478 346 2482
rect 462 2478 466 2482
rect 1406 2478 1410 2482
rect 1590 2478 1594 2482
rect 1614 2478 1618 2482
rect 1678 2478 1682 2482
rect 1686 2478 1690 2482
rect 1742 2478 1746 2482
rect 1806 2478 1810 2482
rect 1822 2478 1826 2482
rect 1862 2478 1866 2482
rect 1902 2478 1906 2482
rect 1942 2478 1946 2482
rect 1990 2478 1994 2482
rect 2046 2478 2050 2482
rect 2070 2478 2074 2482
rect 2078 2478 2082 2482
rect 2110 2478 2114 2482
rect 2254 2478 2258 2482
rect 2342 2478 2346 2482
rect 2406 2478 2410 2482
rect 2454 2478 2458 2482
rect 6 2468 10 2472
rect 54 2468 58 2472
rect 62 2468 66 2472
rect 78 2468 82 2472
rect 94 2468 98 2472
rect 134 2468 138 2472
rect 150 2468 154 2472
rect 182 2468 186 2472
rect 254 2468 258 2472
rect 286 2468 290 2472
rect 302 2468 306 2472
rect 374 2468 378 2472
rect 446 2468 450 2472
rect 494 2468 498 2472
rect 518 2468 522 2472
rect 566 2468 570 2472
rect 598 2468 602 2472
rect 622 2468 626 2472
rect 662 2468 666 2472
rect 742 2468 746 2472
rect 774 2468 778 2472
rect 870 2468 874 2472
rect 878 2468 882 2472
rect 902 2468 906 2472
rect 998 2468 1002 2472
rect 14 2458 18 2462
rect 38 2458 42 2462
rect 102 2458 106 2462
rect 110 2458 114 2462
rect 126 2458 130 2462
rect 174 2458 178 2462
rect 190 2458 194 2462
rect 214 2458 218 2462
rect 270 2458 274 2462
rect 278 2458 282 2462
rect 294 2458 298 2462
rect 326 2458 330 2462
rect 366 2458 370 2462
rect 406 2458 410 2462
rect 414 2458 418 2462
rect 438 2458 442 2462
rect 510 2458 514 2462
rect 574 2458 578 2462
rect 582 2458 586 2462
rect 598 2458 602 2462
rect 670 2458 674 2462
rect 726 2458 730 2462
rect 750 2458 754 2462
rect 766 2458 770 2462
rect 806 2458 810 2462
rect 830 2458 834 2462
rect 838 2458 842 2462
rect 870 2458 874 2462
rect 926 2458 930 2462
rect 934 2458 938 2462
rect 958 2458 962 2462
rect 982 2458 986 2462
rect 990 2458 994 2462
rect 1006 2458 1010 2462
rect 1054 2458 1058 2462
rect 1062 2458 1066 2462
rect 1118 2468 1122 2472
rect 1150 2468 1154 2472
rect 1206 2468 1210 2472
rect 1254 2468 1258 2472
rect 1286 2468 1290 2472
rect 1294 2468 1298 2472
rect 1118 2458 1122 2462
rect 1142 2458 1146 2462
rect 1166 2458 1170 2462
rect 1190 2458 1194 2462
rect 1198 2458 1202 2462
rect 1246 2458 1250 2462
rect 1286 2458 1290 2462
rect 1302 2458 1306 2462
rect 1398 2468 1402 2472
rect 1414 2468 1418 2472
rect 1462 2468 1466 2472
rect 1358 2458 1362 2462
rect 1382 2458 1386 2462
rect 1390 2458 1394 2462
rect 1430 2458 1434 2462
rect 1470 2458 1474 2462
rect 1486 2458 1490 2462
rect 1502 2458 1506 2462
rect 1566 2468 1570 2472
rect 1614 2468 1618 2472
rect 1662 2468 1666 2472
rect 1686 2468 1690 2472
rect 1774 2468 1778 2472
rect 1830 2468 1834 2472
rect 1934 2468 1938 2472
rect 1942 2468 1946 2472
rect 1982 2468 1986 2472
rect 2014 2468 2018 2472
rect 2062 2468 2066 2472
rect 2086 2468 2090 2472
rect 2126 2468 2130 2472
rect 2238 2468 2242 2472
rect 2262 2468 2266 2472
rect 2310 2468 2314 2472
rect 2326 2468 2330 2472
rect 2350 2468 2354 2472
rect 2390 2468 2394 2472
rect 2430 2468 2434 2472
rect 2510 2478 2514 2482
rect 2518 2478 2522 2482
rect 2590 2478 2594 2482
rect 2630 2478 2634 2482
rect 2990 2478 2994 2482
rect 3062 2478 3066 2482
rect 3118 2478 3122 2482
rect 3166 2478 3170 2482
rect 3238 2478 3242 2482
rect 3430 2478 3434 2482
rect 2478 2468 2482 2472
rect 2526 2468 2530 2472
rect 2558 2468 2562 2472
rect 2622 2468 2626 2472
rect 2686 2468 2690 2472
rect 2702 2468 2706 2472
rect 1574 2458 1578 2462
rect 1598 2458 1602 2462
rect 1646 2458 1650 2462
rect 1654 2458 1658 2462
rect 1718 2458 1722 2462
rect 1766 2458 1770 2462
rect 1782 2458 1786 2462
rect 1798 2458 1802 2462
rect 1838 2458 1842 2462
rect 1878 2458 1882 2462
rect 1926 2458 1930 2462
rect 1974 2458 1978 2462
rect 2054 2458 2058 2462
rect 2134 2458 2138 2462
rect 2190 2458 2194 2462
rect 2222 2458 2226 2462
rect 2230 2458 2234 2462
rect 2270 2458 2274 2462
rect 2318 2458 2322 2462
rect 2358 2458 2362 2462
rect 2366 2458 2370 2462
rect 2382 2458 2386 2462
rect 2438 2458 2442 2462
rect 2494 2458 2498 2462
rect 2550 2458 2554 2462
rect 2630 2458 2634 2462
rect 2646 2458 2650 2462
rect 2654 2458 2658 2462
rect 2670 2458 2674 2462
rect 2694 2458 2698 2462
rect 2758 2468 2762 2472
rect 2766 2468 2770 2472
rect 2854 2468 2858 2472
rect 2934 2468 2938 2472
rect 3014 2468 3018 2472
rect 3078 2468 3082 2472
rect 3102 2468 3106 2472
rect 3126 2468 3130 2472
rect 3182 2468 3186 2472
rect 3230 2468 3234 2472
rect 3262 2468 3266 2472
rect 3310 2468 3314 2472
rect 3366 2468 3370 2472
rect 3382 2468 3386 2472
rect 3398 2468 3402 2472
rect 3510 2478 3514 2482
rect 3470 2468 3474 2472
rect 3510 2468 3514 2472
rect 2726 2458 2730 2462
rect 2742 2458 2746 2462
rect 2766 2458 2770 2462
rect 2782 2458 2786 2462
rect 2814 2458 2818 2462
rect 2830 2458 2834 2462
rect 2902 2458 2906 2462
rect 2942 2458 2946 2462
rect 2966 2458 2970 2462
rect 2982 2458 2986 2462
rect 3014 2458 3018 2462
rect 3022 2458 3026 2462
rect 3102 2458 3106 2462
rect 3150 2458 3154 2462
rect 3174 2458 3178 2462
rect 3222 2458 3226 2462
rect 3254 2458 3258 2462
rect 3302 2458 3306 2462
rect 3318 2458 3322 2462
rect 3406 2458 3410 2462
rect 3454 2458 3458 2462
rect 3494 2458 3498 2462
rect 3526 2458 3530 2462
rect 94 2448 98 2452
rect 126 2448 130 2452
rect 158 2448 162 2452
rect 238 2448 242 2452
rect 318 2448 322 2452
rect 422 2448 426 2452
rect 470 2448 474 2452
rect 534 2448 538 2452
rect 542 2448 546 2452
rect 574 2448 578 2452
rect 606 2448 610 2452
rect 686 2448 690 2452
rect 710 2448 714 2452
rect 790 2448 794 2452
rect 846 2448 850 2452
rect 894 2448 898 2452
rect 918 2448 922 2452
rect 974 2448 978 2452
rect 1086 2448 1090 2452
rect 1126 2448 1130 2452
rect 1222 2448 1226 2452
rect 1262 2448 1266 2452
rect 1326 2448 1330 2452
rect 1494 2448 1498 2452
rect 1526 2448 1530 2452
rect 1542 2448 1546 2452
rect 1590 2448 1594 2452
rect 1678 2448 1682 2452
rect 1750 2448 1754 2452
rect 1814 2448 1818 2452
rect 1854 2448 1858 2452
rect 1910 2448 1914 2452
rect 1958 2448 1962 2452
rect 2102 2448 2106 2452
rect 2158 2448 2162 2452
rect 2286 2448 2290 2452
rect 2294 2448 2298 2452
rect 2374 2448 2378 2452
rect 2414 2448 2418 2452
rect 2598 2448 2602 2452
rect 2678 2448 2682 2452
rect 2734 2448 2738 2452
rect 2750 2448 2754 2452
rect 2790 2448 2794 2452
rect 2822 2448 2826 2452
rect 2958 2448 2962 2452
rect 2966 2448 2970 2452
rect 3022 2448 3026 2452
rect 3038 2448 3042 2452
rect 3078 2448 3082 2452
rect 3118 2448 3122 2452
rect 3142 2448 3146 2452
rect 3206 2448 3210 2452
rect 3278 2448 3282 2452
rect 3374 2448 3378 2452
rect 3518 2448 3522 2452
rect 462 2438 466 2442
rect 502 2438 506 2442
rect 1094 2438 1098 2442
rect 1510 2438 1514 2442
rect 1558 2438 1562 2442
rect 1766 2438 1770 2442
rect 2254 2438 2258 2442
rect 2342 2438 2346 2442
rect 2550 2438 2554 2442
rect 2734 2438 2738 2442
rect 2806 2438 2810 2442
rect 3534 2438 3538 2442
rect 1142 2428 1146 2432
rect 1422 2428 1426 2432
rect 14 2418 18 2422
rect 358 2418 362 2422
rect 398 2418 402 2422
rect 438 2418 442 2422
rect 486 2418 490 2422
rect 558 2418 562 2422
rect 614 2418 618 2422
rect 646 2418 650 2422
rect 670 2418 674 2422
rect 694 2418 698 2422
rect 750 2418 754 2422
rect 822 2418 826 2422
rect 862 2418 866 2422
rect 886 2418 890 2422
rect 910 2418 914 2422
rect 950 2418 954 2422
rect 1046 2418 1050 2422
rect 1110 2418 1114 2422
rect 1182 2418 1186 2422
rect 1214 2418 1218 2422
rect 1246 2418 1250 2422
rect 1278 2418 1282 2422
rect 1374 2418 1378 2422
rect 1894 2418 1898 2422
rect 1926 2418 1930 2422
rect 2094 2418 2098 2422
rect 2110 2418 2114 2422
rect 2846 2418 2850 2422
rect 2886 2418 2890 2422
rect 3070 2418 3074 2422
rect 3246 2418 3250 2422
rect 3526 2418 3530 2422
rect 482 2403 486 2407
rect 489 2403 493 2407
rect 1514 2403 1518 2407
rect 1521 2403 1525 2407
rect 2538 2403 2542 2407
rect 2545 2403 2549 2407
rect 918 2388 922 2392
rect 1326 2388 1330 2392
rect 1422 2388 1426 2392
rect 1566 2388 1570 2392
rect 1806 2388 1810 2392
rect 1854 2388 1858 2392
rect 1886 2388 1890 2392
rect 2070 2388 2074 2392
rect 2134 2388 2138 2392
rect 2374 2388 2378 2392
rect 2406 2388 2410 2392
rect 2510 2388 2514 2392
rect 2710 2388 2714 2392
rect 2734 2388 2738 2392
rect 2870 2388 2874 2392
rect 3094 2388 3098 2392
rect 3118 2388 3122 2392
rect 3390 2388 3394 2392
rect 3518 2388 3522 2392
rect 318 2378 322 2382
rect 342 2368 346 2372
rect 406 2368 410 2372
rect 614 2368 618 2372
rect 758 2368 762 2372
rect 1334 2368 1338 2372
rect 2062 2368 2066 2372
rect 2158 2368 2162 2372
rect 2230 2368 2234 2372
rect 2286 2368 2290 2372
rect 2366 2368 2370 2372
rect 2790 2368 2794 2372
rect 2934 2368 2938 2372
rect 3294 2368 3298 2372
rect 6 2358 10 2362
rect 54 2358 58 2362
rect 62 2358 66 2362
rect 118 2358 122 2362
rect 174 2358 178 2362
rect 230 2358 234 2362
rect 238 2358 242 2362
rect 286 2358 290 2362
rect 38 2348 42 2352
rect 78 2348 82 2352
rect 102 2348 106 2352
rect 126 2348 130 2352
rect 134 2348 138 2352
rect 158 2348 162 2352
rect 190 2348 194 2352
rect 214 2348 218 2352
rect 254 2348 258 2352
rect 358 2358 362 2362
rect 366 2358 370 2362
rect 462 2358 466 2362
rect 502 2358 506 2362
rect 542 2358 546 2362
rect 550 2358 554 2362
rect 630 2358 634 2362
rect 638 2358 642 2362
rect 670 2358 674 2362
rect 702 2358 706 2362
rect 734 2358 738 2362
rect 750 2358 754 2362
rect 790 2358 794 2362
rect 846 2358 850 2362
rect 854 2358 858 2362
rect 886 2358 890 2362
rect 998 2358 1002 2362
rect 1030 2358 1034 2362
rect 342 2348 346 2352
rect 406 2348 410 2352
rect 566 2348 570 2352
rect 590 2348 594 2352
rect 654 2348 658 2352
rect 670 2348 674 2352
rect 686 2348 690 2352
rect 718 2348 722 2352
rect 774 2348 778 2352
rect 790 2348 794 2352
rect 806 2348 810 2352
rect 822 2348 826 2352
rect 830 2348 834 2352
rect 870 2348 874 2352
rect 886 2348 890 2352
rect 902 2348 906 2352
rect 942 2348 946 2352
rect 974 2348 978 2352
rect 998 2348 1002 2352
rect 1046 2348 1050 2352
rect 1070 2358 1074 2362
rect 1094 2358 1098 2362
rect 1142 2358 1146 2362
rect 1214 2358 1218 2362
rect 1110 2348 1114 2352
rect 1150 2348 1154 2352
rect 1158 2348 1162 2352
rect 1190 2348 1194 2352
rect 1278 2358 1282 2362
rect 1302 2358 1306 2362
rect 1350 2358 1354 2362
rect 1374 2358 1378 2362
rect 1238 2348 1242 2352
rect 1246 2348 1250 2352
rect 1342 2348 1346 2352
rect 1454 2358 1458 2362
rect 1486 2358 1490 2362
rect 1598 2358 1602 2362
rect 1398 2348 1402 2352
rect 1438 2348 1442 2352
rect 1470 2348 1474 2352
rect 1526 2348 1530 2352
rect 1534 2348 1538 2352
rect 1614 2348 1618 2352
rect 1662 2348 1666 2352
rect 1694 2348 1698 2352
rect 1718 2358 1722 2362
rect 1750 2358 1754 2362
rect 1918 2358 1922 2362
rect 1982 2358 1986 2362
rect 2142 2358 2146 2362
rect 2198 2358 2202 2362
rect 2246 2358 2250 2362
rect 2350 2358 2354 2362
rect 2382 2358 2386 2362
rect 2390 2358 2394 2362
rect 2502 2358 2506 2362
rect 2590 2358 2594 2362
rect 2646 2358 2650 2362
rect 2750 2358 2754 2362
rect 2814 2358 2818 2362
rect 2862 2358 2866 2362
rect 2950 2358 2954 2362
rect 2958 2358 2962 2362
rect 3070 2358 3074 2362
rect 3158 2358 3162 2362
rect 3174 2358 3178 2362
rect 3230 2358 3234 2362
rect 3406 2358 3410 2362
rect 3438 2358 3442 2362
rect 3470 2358 3474 2362
rect 1734 2348 1738 2352
rect 1766 2348 1770 2352
rect 1782 2348 1786 2352
rect 1798 2348 1802 2352
rect 1854 2348 1858 2352
rect 1910 2348 1914 2352
rect 1926 2348 1930 2352
rect 1966 2348 1970 2352
rect 2006 2348 2010 2352
rect 2038 2348 2042 2352
rect 2070 2348 2074 2352
rect 2198 2348 2202 2352
rect 2230 2348 2234 2352
rect 2286 2348 2290 2352
rect 2318 2348 2322 2352
rect 2334 2348 2338 2352
rect 2342 2348 2346 2352
rect 2374 2348 2378 2352
rect 2414 2348 2418 2352
rect 2470 2348 2474 2352
rect 2534 2348 2538 2352
rect 2582 2348 2586 2352
rect 2606 2348 2610 2352
rect 2622 2348 2626 2352
rect 2630 2348 2634 2352
rect 2654 2348 2658 2352
rect 2686 2348 2690 2352
rect 2694 2348 2698 2352
rect 2718 2348 2722 2352
rect 2734 2348 2738 2352
rect 2830 2348 2834 2352
rect 22 2338 26 2342
rect 30 2338 34 2342
rect 86 2338 90 2342
rect 94 2338 98 2342
rect 182 2338 186 2342
rect 198 2338 202 2342
rect 222 2338 226 2342
rect 302 2338 306 2342
rect 334 2338 338 2342
rect 382 2338 386 2342
rect 390 2338 394 2342
rect 414 2338 418 2342
rect 446 2338 450 2342
rect 470 2338 474 2342
rect 526 2338 530 2342
rect 582 2338 586 2342
rect 614 2338 618 2342
rect 662 2338 666 2342
rect 694 2338 698 2342
rect 726 2338 730 2342
rect 734 2338 738 2342
rect 782 2338 786 2342
rect 814 2338 818 2342
rect 894 2338 898 2342
rect 910 2338 914 2342
rect 926 2338 930 2342
rect 934 2338 938 2342
rect 966 2338 970 2342
rect 1014 2338 1018 2342
rect 1038 2338 1042 2342
rect 1054 2338 1058 2342
rect 1086 2338 1090 2342
rect 1102 2338 1106 2342
rect 1118 2338 1122 2342
rect 1126 2338 1130 2342
rect 1190 2338 1194 2342
rect 1254 2338 1258 2342
rect 1286 2338 1290 2342
rect 1302 2338 1306 2342
rect 1358 2338 1362 2342
rect 1406 2338 1410 2342
rect 1462 2338 1466 2342
rect 1502 2338 1506 2342
rect 1550 2338 1554 2342
rect 1574 2338 1578 2342
rect 1598 2338 1602 2342
rect 1614 2338 1618 2342
rect 1654 2338 1658 2342
rect 1710 2338 1714 2342
rect 1742 2338 1746 2342
rect 1774 2338 1778 2342
rect 1822 2338 1826 2342
rect 1862 2338 1866 2342
rect 1942 2338 1946 2342
rect 2102 2338 2106 2342
rect 2110 2338 2114 2342
rect 2134 2338 2138 2342
rect 2158 2338 2162 2342
rect 2182 2338 2186 2342
rect 2214 2338 2218 2342
rect 2222 2338 2226 2342
rect 2270 2338 2274 2342
rect 2318 2338 2322 2342
rect 2414 2338 2418 2342
rect 2422 2338 2426 2342
rect 2470 2338 2474 2342
rect 2478 2338 2482 2342
rect 2494 2338 2498 2342
rect 2574 2338 2578 2342
rect 2622 2338 2626 2342
rect 2662 2338 2666 2342
rect 2678 2338 2682 2342
rect 2726 2338 2730 2342
rect 2758 2338 2762 2342
rect 2806 2338 2810 2342
rect 2822 2338 2826 2342
rect 2838 2338 2842 2342
rect 2886 2338 2890 2342
rect 2902 2348 2906 2352
rect 2934 2348 2938 2352
rect 2958 2348 2962 2352
rect 2982 2348 2986 2352
rect 3094 2348 3098 2352
rect 3158 2348 3162 2352
rect 3182 2348 3186 2352
rect 3214 2348 3218 2352
rect 3254 2348 3258 2352
rect 3326 2348 3330 2352
rect 3342 2348 3346 2352
rect 3350 2348 3354 2352
rect 3382 2348 3386 2352
rect 3414 2348 3418 2352
rect 3454 2348 3458 2352
rect 3478 2348 3482 2352
rect 3510 2348 3514 2352
rect 3526 2348 3530 2352
rect 2926 2338 2930 2342
rect 2998 2338 3002 2342
rect 3038 2338 3042 2342
rect 3102 2338 3106 2342
rect 3110 2338 3114 2342
rect 3142 2338 3146 2342
rect 3158 2338 3162 2342
rect 3174 2338 3178 2342
rect 3206 2338 3210 2342
rect 3262 2338 3266 2342
rect 3310 2338 3314 2342
rect 3334 2338 3338 2342
rect 3358 2338 3362 2342
rect 3366 2338 3370 2342
rect 3382 2338 3386 2342
rect 3422 2338 3426 2342
rect 3438 2338 3442 2342
rect 3558 2338 3562 2342
rect 278 2328 282 2332
rect 478 2328 482 2332
rect 518 2328 522 2332
rect 1454 2328 1458 2332
rect 1518 2328 1522 2332
rect 1566 2328 1570 2332
rect 1630 2328 1634 2332
rect 1654 2328 1658 2332
rect 1678 2328 1682 2332
rect 1750 2328 1754 2332
rect 1782 2328 1786 2332
rect 1830 2328 1834 2332
rect 1838 2328 1842 2332
rect 1862 2328 1866 2332
rect 1894 2328 1898 2332
rect 1910 2328 1914 2332
rect 1950 2328 1954 2332
rect 1966 2328 1970 2332
rect 1982 2328 1986 2332
rect 2006 2328 2010 2332
rect 2030 2328 2034 2332
rect 2118 2328 2122 2332
rect 2166 2328 2170 2332
rect 2318 2328 2322 2332
rect 2510 2328 2514 2332
rect 2558 2328 2562 2332
rect 2590 2328 2594 2332
rect 2662 2328 2666 2332
rect 2870 2328 2874 2332
rect 2918 2328 2922 2332
rect 3006 2328 3010 2332
rect 3054 2328 3058 2332
rect 3126 2328 3130 2332
rect 3222 2328 3226 2332
rect 3238 2328 3242 2332
rect 3318 2328 3322 2332
rect 3374 2328 3378 2332
rect 3438 2328 3442 2332
rect 3526 2328 3530 2332
rect 6 2318 10 2322
rect 54 2318 58 2322
rect 62 2318 66 2322
rect 118 2318 122 2322
rect 150 2318 154 2322
rect 238 2318 242 2322
rect 294 2318 298 2322
rect 374 2318 378 2322
rect 398 2318 402 2322
rect 438 2318 442 2322
rect 510 2318 514 2322
rect 534 2318 538 2322
rect 550 2318 554 2322
rect 606 2318 610 2322
rect 638 2318 642 2322
rect 702 2318 706 2322
rect 758 2318 762 2322
rect 846 2318 850 2322
rect 854 2318 858 2322
rect 918 2318 922 2322
rect 958 2318 962 2322
rect 1030 2318 1034 2322
rect 1142 2318 1146 2322
rect 1174 2318 1178 2322
rect 1222 2318 1226 2322
rect 1278 2318 1282 2322
rect 1302 2318 1306 2322
rect 1318 2318 1322 2322
rect 1382 2318 1386 2322
rect 1590 2318 1594 2322
rect 1998 2318 2002 2322
rect 2206 2318 2210 2322
rect 2262 2318 2266 2322
rect 2302 2318 2306 2322
rect 2454 2318 2458 2322
rect 2646 2318 2650 2322
rect 2710 2318 2714 2322
rect 2862 2318 2866 2322
rect 3046 2318 3050 2322
rect 3134 2318 3138 2322
rect 3246 2318 3250 2322
rect 3494 2318 3498 2322
rect 994 2303 998 2307
rect 1001 2303 1005 2307
rect 2026 2303 2030 2307
rect 2033 2303 2037 2307
rect 3042 2303 3046 2307
rect 3049 2303 3053 2307
rect 46 2288 50 2292
rect 358 2288 362 2292
rect 878 2288 882 2292
rect 1542 2288 1546 2292
rect 1798 2288 1802 2292
rect 1838 2288 1842 2292
rect 1902 2288 1906 2292
rect 2046 2288 2050 2292
rect 2078 2288 2082 2292
rect 2118 2288 2122 2292
rect 2150 2288 2154 2292
rect 2358 2288 2362 2292
rect 2566 2288 2570 2292
rect 2590 2288 2594 2292
rect 2646 2288 2650 2292
rect 2782 2288 2786 2292
rect 2918 2288 2922 2292
rect 3030 2288 3034 2292
rect 3150 2288 3154 2292
rect 3174 2288 3178 2292
rect 3310 2288 3314 2292
rect 3334 2288 3338 2292
rect 3390 2288 3394 2292
rect 3550 2288 3554 2292
rect 326 2278 330 2282
rect 30 2268 34 2272
rect 38 2268 42 2272
rect 86 2268 90 2272
rect 286 2268 290 2272
rect 310 2268 314 2272
rect 30 2258 34 2262
rect 94 2258 98 2262
rect 102 2258 106 2262
rect 126 2258 130 2262
rect 134 2258 138 2262
rect 150 2258 154 2262
rect 174 2258 178 2262
rect 182 2258 186 2262
rect 198 2258 202 2262
rect 222 2258 226 2262
rect 230 2258 234 2262
rect 246 2258 250 2262
rect 270 2258 274 2262
rect 278 2258 282 2262
rect 302 2258 306 2262
rect 342 2268 346 2272
rect 358 2268 362 2272
rect 390 2268 394 2272
rect 414 2268 418 2272
rect 382 2258 386 2262
rect 566 2278 570 2282
rect 590 2278 594 2282
rect 606 2278 610 2282
rect 670 2278 674 2282
rect 766 2278 770 2282
rect 790 2278 794 2282
rect 806 2278 810 2282
rect 1454 2278 1458 2282
rect 1470 2278 1474 2282
rect 1478 2278 1482 2282
rect 1494 2278 1498 2282
rect 1510 2278 1514 2282
rect 1534 2278 1538 2282
rect 1614 2278 1618 2282
rect 1806 2278 1810 2282
rect 1814 2278 1818 2282
rect 1846 2278 1850 2282
rect 1894 2278 1898 2282
rect 1966 2278 1970 2282
rect 1982 2278 1986 2282
rect 2158 2278 2162 2282
rect 2198 2278 2202 2282
rect 2222 2278 2226 2282
rect 2334 2278 2338 2282
rect 2366 2278 2370 2282
rect 2382 2278 2386 2282
rect 2598 2278 2602 2282
rect 2678 2278 2682 2282
rect 2798 2278 2802 2282
rect 3350 2278 3354 2282
rect 3398 2278 3402 2282
rect 3486 2278 3490 2282
rect 438 2268 442 2272
rect 462 2268 466 2272
rect 558 2268 562 2272
rect 574 2268 578 2272
rect 678 2268 682 2272
rect 710 2268 714 2272
rect 758 2268 762 2272
rect 782 2268 786 2272
rect 862 2268 866 2272
rect 886 2268 890 2272
rect 910 2268 914 2272
rect 1054 2268 1058 2272
rect 438 2258 442 2262
rect 462 2258 466 2262
rect 494 2258 498 2262
rect 518 2258 522 2262
rect 526 2258 530 2262
rect 550 2258 554 2262
rect 614 2258 618 2262
rect 622 2258 626 2262
rect 646 2258 650 2262
rect 686 2258 690 2262
rect 750 2258 754 2262
rect 822 2258 826 2262
rect 846 2258 850 2262
rect 854 2258 858 2262
rect 902 2258 906 2262
rect 918 2258 922 2262
rect 926 2258 930 2262
rect 950 2258 954 2262
rect 974 2258 978 2262
rect 998 2258 1002 2262
rect 1006 2258 1010 2262
rect 1014 2258 1018 2262
rect 1046 2258 1050 2262
rect 1070 2258 1074 2262
rect 1078 2258 1082 2262
rect 1094 2268 1098 2272
rect 1142 2268 1146 2272
rect 1182 2268 1186 2272
rect 1238 2268 1242 2272
rect 1262 2268 1266 2272
rect 1270 2268 1274 2272
rect 1350 2268 1354 2272
rect 1398 2268 1402 2272
rect 1566 2268 1570 2272
rect 1574 2268 1578 2272
rect 1590 2268 1594 2272
rect 1606 2268 1610 2272
rect 1630 2268 1634 2272
rect 1646 2268 1650 2272
rect 1678 2268 1682 2272
rect 1702 2268 1706 2272
rect 1718 2268 1722 2272
rect 1726 2268 1730 2272
rect 1742 2268 1746 2272
rect 1750 2268 1754 2272
rect 1782 2268 1786 2272
rect 1830 2268 1834 2272
rect 1878 2268 1882 2272
rect 1910 2268 1914 2272
rect 1958 2268 1962 2272
rect 1998 2268 2002 2272
rect 2014 2268 2018 2272
rect 2070 2268 2074 2272
rect 2102 2268 2106 2272
rect 2126 2268 2130 2272
rect 2142 2268 2146 2272
rect 2166 2268 2170 2272
rect 2182 2268 2186 2272
rect 2230 2268 2234 2272
rect 2254 2268 2258 2272
rect 1094 2258 1098 2262
rect 1126 2258 1130 2262
rect 1142 2258 1146 2262
rect 1166 2258 1170 2262
rect 1174 2258 1178 2262
rect 1230 2258 1234 2262
rect 1278 2258 1282 2262
rect 1294 2258 1298 2262
rect 1334 2258 1338 2262
rect 1342 2258 1346 2262
rect 1382 2258 1386 2262
rect 1390 2258 1394 2262
rect 1414 2258 1418 2262
rect 1438 2258 1442 2262
rect 1446 2258 1450 2262
rect 1478 2258 1482 2262
rect 1550 2258 1554 2262
rect 1582 2258 1586 2262
rect 1598 2258 1602 2262
rect 1646 2258 1650 2262
rect 1822 2258 1826 2262
rect 1854 2258 1858 2262
rect 1886 2258 1890 2262
rect 2262 2266 2266 2270
rect 2286 2268 2290 2272
rect 2390 2268 2394 2272
rect 2406 2268 2410 2272
rect 2422 2268 2426 2272
rect 2438 2268 2442 2272
rect 2454 2268 2458 2272
rect 2582 2268 2586 2272
rect 2630 2268 2634 2272
rect 2686 2268 2690 2272
rect 2702 2268 2706 2272
rect 2734 2268 2738 2272
rect 2766 2268 2770 2272
rect 2814 2268 2818 2272
rect 2846 2268 2850 2272
rect 2854 2268 2858 2272
rect 2910 2268 2914 2272
rect 2942 2268 2946 2272
rect 2950 2268 2954 2272
rect 2998 2268 3002 2272
rect 3006 2268 3010 2272
rect 3054 2268 3058 2272
rect 1990 2258 1994 2262
rect 2022 2258 2026 2262
rect 2062 2258 2066 2262
rect 2134 2258 2138 2262
rect 2198 2258 2202 2262
rect 2278 2258 2282 2262
rect 2310 2258 2314 2262
rect 2318 2258 2322 2262
rect 2342 2258 2346 2262
rect 2398 2258 2402 2262
rect 2430 2258 2434 2262
rect 2494 2258 2498 2262
rect 2518 2258 2522 2262
rect 2574 2258 2578 2262
rect 2606 2258 2610 2262
rect 2662 2258 2666 2262
rect 2694 2258 2698 2262
rect 2710 2258 2714 2262
rect 2734 2258 2738 2262
rect 2758 2258 2762 2262
rect 2814 2258 2818 2262
rect 2838 2258 2842 2262
rect 2862 2258 2866 2262
rect 2902 2258 2906 2262
rect 2934 2258 2938 2262
rect 2998 2258 3002 2262
rect 3062 2258 3066 2262
rect 3102 2258 3106 2262
rect 3118 2268 3122 2272
rect 3134 2268 3138 2272
rect 3158 2268 3162 2272
rect 3182 2268 3186 2272
rect 3214 2268 3218 2272
rect 3246 2268 3250 2272
rect 3262 2268 3266 2272
rect 3302 2268 3306 2272
rect 3342 2268 3346 2272
rect 3430 2268 3434 2272
rect 3134 2258 3138 2262
rect 3190 2258 3194 2262
rect 3214 2258 3218 2262
rect 3286 2258 3290 2262
rect 3374 2258 3378 2262
rect 3454 2258 3458 2262
rect 3494 2258 3498 2262
rect 3510 2258 3514 2262
rect 6 2248 10 2252
rect 334 2248 338 2252
rect 358 2248 362 2252
rect 366 2248 370 2252
rect 398 2248 402 2252
rect 430 2248 434 2252
rect 534 2248 538 2252
rect 590 2248 594 2252
rect 878 2248 882 2252
rect 1030 2248 1034 2252
rect 1062 2248 1066 2252
rect 1118 2248 1122 2252
rect 1150 2248 1154 2252
rect 1206 2248 1210 2252
rect 1214 2248 1218 2252
rect 1246 2248 1250 2252
rect 1294 2248 1298 2252
rect 1366 2248 1370 2252
rect 1558 2248 1562 2252
rect 1662 2248 1666 2252
rect 1702 2248 1706 2252
rect 1742 2248 1746 2252
rect 1774 2248 1778 2252
rect 1798 2248 1802 2252
rect 2046 2248 2050 2252
rect 2078 2248 2082 2252
rect 2110 2248 2114 2252
rect 2438 2248 2442 2252
rect 2638 2248 2642 2252
rect 2710 2248 2714 2252
rect 2718 2248 2722 2252
rect 2742 2248 2746 2252
rect 2774 2248 2778 2252
rect 2822 2248 2826 2252
rect 2886 2248 2890 2252
rect 2918 2248 2922 2252
rect 3030 2248 3034 2252
rect 3062 2248 3066 2252
rect 3086 2248 3090 2252
rect 3150 2248 3154 2252
rect 3174 2248 3178 2252
rect 3206 2248 3210 2252
rect 3238 2248 3242 2252
rect 3262 2248 3266 2252
rect 3318 2248 3322 2252
rect 3390 2248 3394 2252
rect 3430 2248 3434 2252
rect 3454 2248 3458 2252
rect 54 2238 58 2242
rect 670 2238 674 2242
rect 686 2238 690 2242
rect 726 2238 730 2242
rect 1942 2238 1946 2242
rect 2206 2238 2210 2242
rect 2254 2238 2258 2242
rect 3222 2238 3226 2242
rect 1254 2228 1258 2232
rect 3422 2228 3426 2232
rect 22 2218 26 2222
rect 78 2218 82 2222
rect 110 2218 114 2222
rect 166 2218 170 2222
rect 206 2218 210 2222
rect 262 2218 266 2222
rect 406 2218 410 2222
rect 422 2218 426 2222
rect 502 2218 506 2222
rect 550 2218 554 2222
rect 582 2218 586 2222
rect 630 2218 634 2222
rect 750 2218 754 2222
rect 774 2218 778 2222
rect 798 2218 802 2222
rect 838 2218 842 2222
rect 942 2218 946 2222
rect 990 2218 994 2222
rect 1166 2218 1170 2222
rect 1190 2218 1194 2222
rect 1230 2218 1234 2222
rect 1278 2218 1282 2222
rect 1326 2218 1330 2222
rect 1422 2218 1426 2222
rect 1614 2218 1618 2222
rect 1758 2218 1762 2222
rect 1878 2218 1882 2222
rect 2014 2218 2018 2222
rect 2422 2218 2426 2222
rect 2558 2218 2562 2222
rect 2862 2218 2866 2222
rect 2966 2218 2970 2222
rect 3190 2218 3194 2222
rect 482 2203 486 2207
rect 489 2203 493 2207
rect 1514 2203 1518 2207
rect 1521 2203 1525 2207
rect 2538 2203 2542 2207
rect 2545 2203 2549 2207
rect 230 2188 234 2192
rect 1766 2188 1770 2192
rect 1894 2188 1898 2192
rect 1966 2188 1970 2192
rect 2046 2188 2050 2192
rect 2270 2188 2274 2192
rect 2334 2188 2338 2192
rect 2486 2188 2490 2192
rect 2574 2188 2578 2192
rect 2758 2188 2762 2192
rect 2798 2188 2802 2192
rect 2974 2188 2978 2192
rect 3182 2188 3186 2192
rect 3270 2188 3274 2192
rect 3390 2188 3394 2192
rect 3470 2188 3474 2192
rect 3542 2188 3546 2192
rect 1518 2178 1522 2182
rect 1718 2178 1722 2182
rect 3102 2178 3106 2182
rect 1534 2168 1538 2172
rect 2126 2168 2130 2172
rect 2150 2168 2154 2172
rect 3150 2168 3154 2172
rect 70 2158 74 2162
rect 110 2158 114 2162
rect 118 2158 122 2162
rect 150 2158 154 2162
rect 190 2158 194 2162
rect 214 2158 218 2162
rect 270 2158 274 2162
rect 278 2158 282 2162
rect 334 2158 338 2162
rect 342 2158 346 2162
rect 366 2158 370 2162
rect 390 2158 394 2162
rect 406 2158 410 2162
rect 6 2148 10 2152
rect 30 2148 34 2152
rect 54 2148 58 2152
rect 62 2148 66 2152
rect 86 2148 90 2152
rect 246 2148 250 2152
rect 302 2148 306 2152
rect 318 2148 322 2152
rect 390 2148 394 2152
rect 430 2148 434 2152
rect 454 2148 458 2152
rect 478 2158 482 2162
rect 542 2158 546 2162
rect 598 2158 602 2162
rect 646 2158 650 2162
rect 678 2158 682 2162
rect 718 2158 722 2162
rect 774 2158 778 2162
rect 822 2158 826 2162
rect 854 2158 858 2162
rect 894 2158 898 2162
rect 958 2158 962 2162
rect 982 2158 986 2162
rect 1054 2158 1058 2162
rect 1078 2158 1082 2162
rect 1134 2158 1138 2162
rect 590 2148 594 2152
rect 630 2148 634 2152
rect 950 2148 954 2152
rect 1190 2158 1194 2162
rect 1254 2158 1258 2162
rect 1262 2158 1266 2162
rect 1286 2158 1290 2162
rect 1310 2158 1314 2162
rect 1350 2158 1354 2162
rect 1374 2158 1378 2162
rect 1158 2148 1162 2152
rect 1166 2148 1170 2152
rect 1198 2148 1202 2152
rect 1222 2148 1226 2152
rect 1286 2148 1290 2152
rect 1414 2158 1418 2162
rect 1550 2158 1554 2162
rect 1598 2158 1602 2162
rect 1606 2158 1610 2162
rect 1638 2158 1642 2162
rect 1670 2158 1674 2162
rect 1750 2158 1754 2162
rect 1878 2158 1882 2162
rect 1910 2158 1914 2162
rect 1982 2158 1986 2162
rect 2006 2158 2010 2162
rect 2110 2158 2114 2162
rect 2222 2158 2226 2162
rect 2254 2158 2258 2162
rect 2350 2158 2354 2162
rect 2406 2158 2410 2162
rect 2518 2158 2522 2162
rect 2726 2158 2730 2162
rect 2806 2158 2810 2162
rect 2822 2158 2826 2162
rect 2838 2158 2842 2162
rect 2910 2158 2914 2162
rect 2918 2158 2922 2162
rect 2934 2158 2938 2162
rect 2958 2158 2962 2162
rect 1438 2148 1442 2152
rect 1446 2148 1450 2152
rect 1470 2148 1474 2152
rect 1486 2148 1490 2152
rect 1518 2148 1522 2152
rect 1534 2148 1538 2152
rect 1558 2148 1562 2152
rect 1622 2148 1626 2152
rect 1654 2148 1658 2152
rect 1782 2148 1786 2152
rect 1798 2148 1802 2152
rect 1830 2148 1834 2152
rect 1862 2148 1866 2152
rect 1894 2148 1898 2152
rect 1910 2148 1914 2152
rect 1966 2148 1970 2152
rect 2030 2148 2034 2152
rect 86 2138 90 2142
rect 94 2138 98 2142
rect 150 2138 154 2142
rect 166 2138 170 2142
rect 174 2138 178 2142
rect 198 2138 202 2142
rect 254 2138 258 2142
rect 310 2138 314 2142
rect 326 2138 330 2142
rect 358 2138 362 2142
rect 390 2138 394 2142
rect 406 2138 410 2142
rect 446 2138 450 2142
rect 518 2138 522 2142
rect 566 2138 570 2142
rect 614 2138 618 2142
rect 622 2138 626 2142
rect 638 2138 642 2142
rect 654 2138 658 2142
rect 694 2138 698 2142
rect 702 2138 706 2142
rect 726 2138 730 2142
rect 758 2138 762 2142
rect 798 2138 802 2142
rect 806 2138 810 2142
rect 830 2138 834 2142
rect 870 2138 874 2142
rect 878 2138 882 2142
rect 918 2138 922 2142
rect 926 2138 930 2142
rect 974 2138 978 2142
rect 998 2138 1002 2142
rect 1046 2138 1050 2142
rect 1070 2138 1074 2142
rect 1094 2138 1098 2142
rect 1118 2138 1122 2142
rect 1174 2138 1178 2142
rect 1222 2138 1226 2142
rect 1246 2138 1250 2142
rect 1278 2138 1282 2142
rect 1302 2138 1306 2142
rect 1326 2138 1330 2142
rect 1334 2138 1338 2142
rect 1358 2138 1362 2142
rect 1382 2138 1386 2142
rect 1430 2138 1434 2142
rect 1582 2138 1586 2142
rect 1630 2138 1634 2142
rect 1646 2138 1650 2142
rect 1670 2138 1674 2142
rect 1694 2138 1698 2142
rect 1734 2138 1738 2142
rect 1790 2138 1794 2142
rect 1822 2138 1826 2142
rect 1854 2138 1858 2142
rect 1886 2138 1890 2142
rect 1950 2138 1954 2142
rect 1958 2138 1962 2142
rect 1990 2138 1994 2142
rect 2006 2138 2010 2142
rect 2070 2138 2074 2142
rect 2086 2148 2090 2152
rect 2126 2148 2130 2152
rect 2142 2148 2146 2152
rect 2174 2148 2178 2152
rect 2190 2148 2194 2152
rect 2206 2148 2210 2152
rect 2238 2148 2242 2152
rect 2278 2148 2282 2152
rect 2286 2148 2290 2152
rect 2302 2148 2306 2152
rect 2318 2148 2322 2152
rect 2366 2148 2370 2152
rect 2390 2148 2394 2152
rect 2414 2148 2418 2152
rect 2430 2148 2434 2152
rect 2462 2148 2466 2152
rect 2502 2148 2506 2152
rect 2558 2148 2562 2152
rect 2598 2148 2602 2152
rect 2622 2148 2626 2152
rect 2630 2148 2634 2152
rect 2662 2148 2666 2152
rect 2694 2148 2698 2152
rect 2702 2148 2706 2152
rect 2742 2148 2746 2152
rect 2774 2148 2778 2152
rect 2822 2148 2826 2152
rect 2854 2148 2858 2152
rect 2870 2148 2874 2152
rect 2886 2148 2890 2152
rect 2918 2148 2922 2152
rect 2934 2148 2938 2152
rect 2942 2148 2946 2152
rect 2990 2158 2994 2162
rect 3014 2158 3018 2162
rect 3070 2158 3074 2162
rect 3166 2158 3170 2162
rect 3206 2158 3210 2162
rect 3238 2158 3242 2162
rect 3286 2158 3290 2162
rect 3326 2158 3330 2162
rect 3406 2158 3410 2162
rect 3070 2148 3074 2152
rect 3158 2148 3162 2152
rect 3198 2148 3202 2152
rect 3222 2148 3226 2152
rect 3254 2148 3258 2152
rect 3342 2148 3346 2152
rect 3358 2148 3362 2152
rect 3390 2148 3394 2152
rect 3414 2148 3418 2152
rect 3430 2148 3434 2152
rect 2166 2138 2170 2142
rect 2198 2138 2202 2142
rect 2230 2138 2234 2142
rect 2310 2138 2314 2142
rect 2326 2138 2330 2142
rect 2374 2138 2378 2142
rect 2494 2138 2498 2142
rect 2606 2138 2610 2142
rect 2670 2138 2674 2142
rect 2686 2138 2690 2142
rect 2694 2138 2698 2142
rect 2742 2138 2746 2142
rect 2766 2138 2770 2142
rect 2782 2138 2786 2142
rect 2830 2138 2834 2142
rect 2862 2138 2866 2142
rect 2894 2138 2898 2142
rect 2942 2138 2946 2142
rect 2966 2138 2970 2142
rect 2998 2138 3002 2142
rect 3030 2138 3034 2142
rect 3078 2138 3082 2142
rect 3086 2138 3090 2142
rect 3134 2138 3138 2142
rect 3230 2138 3234 2142
rect 3254 2138 3258 2142
rect 3262 2138 3266 2142
rect 3310 2138 3314 2142
rect 3350 2138 3354 2142
rect 3382 2138 3386 2142
rect 3422 2138 3426 2142
rect 3438 2138 3442 2142
rect 3478 2138 3482 2142
rect 3486 2138 3490 2142
rect 6 2128 10 2132
rect 158 2128 162 2132
rect 342 2128 346 2132
rect 1110 2128 1114 2132
rect 1510 2128 1514 2132
rect 1574 2128 1578 2132
rect 1918 2128 1922 2132
rect 2102 2128 2106 2132
rect 2262 2128 2266 2132
rect 2414 2128 2418 2132
rect 2430 2128 2434 2132
rect 2454 2128 2458 2132
rect 2486 2128 2490 2132
rect 2526 2128 2530 2132
rect 2718 2128 2722 2132
rect 2798 2128 2802 2132
rect 2870 2128 2874 2132
rect 2958 2128 2962 2132
rect 3294 2128 3298 2132
rect 3374 2128 3378 2132
rect 3462 2128 3466 2132
rect 38 2118 42 2122
rect 110 2118 114 2122
rect 118 2118 122 2122
rect 190 2118 194 2122
rect 206 2118 210 2122
rect 262 2118 266 2122
rect 278 2118 282 2122
rect 366 2118 370 2122
rect 414 2118 418 2122
rect 470 2118 474 2122
rect 534 2118 538 2122
rect 542 2118 546 2122
rect 574 2118 578 2122
rect 598 2118 602 2122
rect 662 2118 666 2122
rect 678 2118 682 2122
rect 718 2118 722 2122
rect 750 2118 754 2122
rect 782 2118 786 2122
rect 822 2118 826 2122
rect 838 2118 842 2122
rect 854 2118 858 2122
rect 886 2118 890 2122
rect 910 2118 914 2122
rect 958 2118 962 2122
rect 1014 2118 1018 2122
rect 1054 2118 1058 2122
rect 1078 2118 1082 2122
rect 1102 2118 1106 2122
rect 1142 2118 1146 2122
rect 1190 2118 1194 2122
rect 1262 2118 1266 2122
rect 1310 2118 1314 2122
rect 1350 2118 1354 2122
rect 1374 2118 1378 2122
rect 1406 2118 1410 2122
rect 1462 2118 1466 2122
rect 1566 2118 1570 2122
rect 1606 2118 1610 2122
rect 1678 2118 1682 2122
rect 1742 2118 1746 2122
rect 1814 2118 1818 2122
rect 1846 2118 1850 2122
rect 1878 2118 1882 2122
rect 1942 2118 1946 2122
rect 2006 2118 2010 2122
rect 2222 2118 2226 2122
rect 2254 2118 2258 2122
rect 2334 2118 2338 2122
rect 2350 2118 2354 2122
rect 2518 2118 2522 2122
rect 2534 2118 2538 2122
rect 2646 2118 2650 2122
rect 2678 2118 2682 2122
rect 2838 2118 2842 2122
rect 3142 2118 3146 2122
rect 3182 2118 3186 2122
rect 3206 2118 3210 2122
rect 3238 2118 3242 2122
rect 3302 2118 3306 2122
rect 3366 2118 3370 2122
rect 3542 2118 3546 2122
rect 994 2103 998 2107
rect 1001 2103 1005 2107
rect 2026 2103 2030 2107
rect 2033 2103 2037 2107
rect 3042 2103 3046 2107
rect 3049 2103 3053 2107
rect 1438 2088 1442 2092
rect 1790 2088 1794 2092
rect 1862 2088 1866 2092
rect 1926 2088 1930 2092
rect 1958 2088 1962 2092
rect 2014 2088 2018 2092
rect 2174 2088 2178 2092
rect 2214 2088 2218 2092
rect 2238 2088 2242 2092
rect 2278 2088 2282 2092
rect 2502 2088 2506 2092
rect 2606 2088 2610 2092
rect 2630 2088 2634 2092
rect 2718 2088 2722 2092
rect 2726 2088 2730 2092
rect 2830 2088 2834 2092
rect 3166 2088 3170 2092
rect 3214 2088 3218 2092
rect 126 2078 130 2082
rect 238 2078 242 2082
rect 286 2078 290 2082
rect 302 2078 306 2082
rect 558 2078 562 2082
rect 790 2078 794 2082
rect 838 2078 842 2082
rect 918 2078 922 2082
rect 1102 2078 1106 2082
rect 1342 2078 1346 2082
rect 1446 2078 1450 2082
rect 1630 2078 1634 2082
rect 1686 2078 1690 2082
rect 1806 2078 1810 2082
rect 1854 2078 1858 2082
rect 1918 2078 1922 2082
rect 1974 2078 1978 2082
rect 6 2068 10 2072
rect 54 2068 58 2072
rect 46 2058 50 2062
rect 86 2068 90 2072
rect 158 2068 162 2072
rect 166 2068 170 2072
rect 270 2068 274 2072
rect 310 2068 314 2072
rect 342 2068 346 2072
rect 438 2068 442 2072
rect 446 2068 450 2072
rect 470 2068 474 2072
rect 494 2068 498 2072
rect 518 2068 522 2072
rect 590 2068 594 2072
rect 646 2068 650 2072
rect 670 2068 674 2072
rect 694 2068 698 2072
rect 758 2068 762 2072
rect 902 2068 906 2072
rect 950 2068 954 2072
rect 982 2068 986 2072
rect 1006 2068 1010 2072
rect 1038 2068 1042 2072
rect 1086 2068 1090 2072
rect 1110 2068 1114 2072
rect 1142 2068 1146 2072
rect 1166 2068 1170 2072
rect 1222 2068 1226 2072
rect 1262 2068 1266 2072
rect 1286 2068 1290 2072
rect 1310 2068 1314 2072
rect 1334 2068 1338 2072
rect 1454 2068 1458 2072
rect 1486 2068 1490 2072
rect 1590 2068 1594 2072
rect 1622 2068 1626 2072
rect 1638 2068 1642 2072
rect 1662 2068 1666 2072
rect 1718 2068 1722 2072
rect 1774 2068 1778 2072
rect 1822 2068 1826 2072
rect 1878 2068 1882 2072
rect 1934 2068 1938 2072
rect 1950 2068 1954 2072
rect 1982 2068 1986 2072
rect 2022 2068 2026 2072
rect 2062 2078 2066 2082
rect 2166 2078 2170 2082
rect 2206 2078 2210 2082
rect 2286 2078 2290 2082
rect 2302 2078 2306 2082
rect 2414 2078 2418 2082
rect 2446 2078 2450 2082
rect 2510 2078 2514 2082
rect 2542 2078 2546 2082
rect 2550 2078 2554 2082
rect 2766 2078 2770 2082
rect 2814 2078 2818 2082
rect 2062 2068 2066 2072
rect 2070 2068 2074 2072
rect 2102 2068 2106 2072
rect 2118 2068 2122 2072
rect 2222 2068 2226 2072
rect 2230 2068 2234 2072
rect 2294 2068 2298 2072
rect 2326 2068 2330 2072
rect 2334 2068 2338 2072
rect 2382 2068 2386 2072
rect 2398 2068 2402 2072
rect 2430 2068 2434 2072
rect 2454 2068 2458 2072
rect 2486 2068 2490 2072
rect 2534 2068 2538 2072
rect 2614 2068 2618 2072
rect 2670 2068 2674 2072
rect 2678 2068 2682 2072
rect 2734 2068 2738 2072
rect 2758 2068 2762 2072
rect 2782 2068 2786 2072
rect 2854 2078 2858 2082
rect 2910 2078 2914 2082
rect 3078 2078 3082 2082
rect 3230 2078 3234 2082
rect 3246 2078 3250 2082
rect 3262 2078 3266 2082
rect 3398 2078 3402 2082
rect 3518 2078 3522 2082
rect 2886 2068 2890 2072
rect 2902 2068 2906 2072
rect 2926 2068 2930 2072
rect 2966 2068 2970 2072
rect 3030 2068 3034 2072
rect 3054 2068 3058 2072
rect 3078 2068 3082 2072
rect 3102 2068 3106 2072
rect 3150 2068 3154 2072
rect 3198 2068 3202 2072
rect 3222 2068 3226 2072
rect 3270 2068 3274 2072
rect 3318 2068 3322 2072
rect 3382 2068 3386 2072
rect 3446 2068 3450 2072
rect 94 2058 98 2062
rect 142 2058 146 2062
rect 150 2058 154 2062
rect 174 2058 178 2062
rect 198 2058 202 2062
rect 214 2058 218 2062
rect 262 2058 266 2062
rect 318 2058 322 2062
rect 350 2058 354 2062
rect 358 2058 362 2062
rect 374 2058 378 2062
rect 382 2058 386 2062
rect 406 2058 410 2062
rect 454 2058 458 2062
rect 526 2058 530 2062
rect 574 2058 578 2062
rect 590 2058 594 2062
rect 598 2058 602 2062
rect 606 2058 610 2062
rect 630 2058 634 2062
rect 646 2058 650 2062
rect 710 2058 714 2062
rect 718 2058 722 2062
rect 734 2058 738 2062
rect 766 2058 770 2062
rect 806 2058 810 2062
rect 862 2058 866 2062
rect 942 2058 946 2062
rect 950 2058 954 2062
rect 974 2058 978 2062
rect 1046 2058 1050 2062
rect 1118 2058 1122 2062
rect 1134 2058 1138 2062
rect 1174 2058 1178 2062
rect 1214 2058 1218 2062
rect 1222 2058 1226 2062
rect 1246 2058 1250 2062
rect 1326 2058 1330 2062
rect 1366 2058 1370 2062
rect 1390 2058 1394 2062
rect 1398 2058 1402 2062
rect 1422 2058 1426 2062
rect 1446 2058 1450 2062
rect 1462 2058 1466 2062
rect 1502 2058 1506 2062
rect 1534 2058 1538 2062
rect 1566 2058 1570 2062
rect 1614 2058 1618 2062
rect 1702 2058 1706 2062
rect 1726 2058 1730 2062
rect 1758 2058 1762 2062
rect 1774 2058 1778 2062
rect 1830 2058 1834 2062
rect 1838 2058 1842 2062
rect 1894 2058 1898 2062
rect 1910 2058 1914 2062
rect 1942 2058 1946 2062
rect 2094 2058 2098 2062
rect 2126 2058 2130 2062
rect 2142 2058 2146 2062
rect 2182 2058 2186 2062
rect 2190 2058 2194 2062
rect 2270 2058 2274 2062
rect 2302 2058 2306 2062
rect 2318 2058 2322 2062
rect 2390 2058 2394 2062
rect 2422 2058 2426 2062
rect 2462 2058 2466 2062
rect 2646 2058 2650 2062
rect 2670 2058 2674 2062
rect 2790 2058 2794 2062
rect 2798 2058 2802 2062
rect 2846 2058 2850 2062
rect 2870 2058 2874 2062
rect 2894 2058 2898 2062
rect 2918 2058 2922 2062
rect 2934 2058 2938 2062
rect 2958 2058 2962 2062
rect 2998 2058 3002 2062
rect 3022 2058 3026 2062
rect 3046 2058 3050 2062
rect 3070 2058 3074 2062
rect 3094 2058 3098 2062
rect 3134 2058 3138 2062
rect 3326 2058 3330 2062
rect 3350 2058 3354 2062
rect 3358 2058 3362 2062
rect 3430 2059 3434 2063
rect 3462 2058 3466 2062
rect 3502 2058 3506 2062
rect 3526 2058 3530 2062
rect 22 2048 26 2052
rect 78 2048 82 2052
rect 110 2048 114 2052
rect 134 2048 138 2052
rect 190 2048 194 2052
rect 198 2048 202 2052
rect 246 2048 250 2052
rect 334 2048 338 2052
rect 366 2048 370 2052
rect 478 2048 482 2052
rect 542 2048 546 2052
rect 566 2048 570 2052
rect 662 2048 666 2052
rect 686 2048 690 2052
rect 750 2048 754 2052
rect 782 2048 786 2052
rect 830 2048 834 2052
rect 886 2048 890 2052
rect 926 2048 930 2052
rect 958 2048 962 2052
rect 1030 2048 1034 2052
rect 1070 2048 1074 2052
rect 1190 2048 1194 2052
rect 1198 2048 1202 2052
rect 1230 2048 1234 2052
rect 1278 2048 1282 2052
rect 1302 2048 1306 2052
rect 1382 2048 1386 2052
rect 1502 2048 1506 2052
rect 1574 2048 1578 2052
rect 1678 2048 1682 2052
rect 1742 2048 1746 2052
rect 1782 2048 1786 2052
rect 1878 2048 1882 2052
rect 1966 2048 1970 2052
rect 2006 2048 2010 2052
rect 2134 2048 2138 2052
rect 2414 2048 2418 2052
rect 2478 2048 2482 2052
rect 2654 2048 2658 2052
rect 2702 2048 2706 2052
rect 2718 2048 2722 2052
rect 2742 2048 2746 2052
rect 2878 2048 2882 2052
rect 2942 2048 2946 2052
rect 2974 2048 2978 2052
rect 2990 2048 2994 2052
rect 3006 2048 3010 2052
rect 3110 2048 3114 2052
rect 3142 2048 3146 2052
rect 3206 2048 3210 2052
rect 3358 2048 3362 2052
rect 1014 2038 1018 2042
rect 1414 2038 1418 2042
rect 1862 2038 1866 2042
rect 1902 2038 1906 2042
rect 2118 2038 2122 2042
rect 2150 2038 2154 2042
rect 2366 2038 2370 2042
rect 2446 2038 2450 2042
rect 2590 2038 2594 2042
rect 2750 2038 2754 2042
rect 2758 2038 2762 2042
rect 3126 2038 3130 2042
rect 3182 2038 3186 2042
rect 3286 2038 3290 2042
rect 3558 2038 3562 2042
rect 46 2018 50 2022
rect 70 2018 74 2022
rect 94 2018 98 2022
rect 118 2018 122 2022
rect 174 2018 178 2022
rect 262 2018 266 2022
rect 278 2018 282 2022
rect 294 2018 298 2022
rect 318 2018 322 2022
rect 398 2018 402 2022
rect 430 2018 434 2022
rect 526 2018 530 2022
rect 550 2018 554 2022
rect 622 2018 626 2022
rect 654 2018 658 2022
rect 734 2018 738 2022
rect 766 2018 770 2022
rect 814 2018 818 2022
rect 862 2018 866 2022
rect 910 2018 914 2022
rect 942 2018 946 2022
rect 1046 2018 1050 2022
rect 1094 2018 1098 2022
rect 1174 2018 1178 2022
rect 1214 2018 1218 2022
rect 1270 2018 1274 2022
rect 1366 2018 1370 2022
rect 1462 2018 1466 2022
rect 1542 2018 1546 2022
rect 1614 2018 1618 2022
rect 1654 2018 1658 2022
rect 1726 2018 1730 2022
rect 1846 2018 1850 2022
rect 1998 2018 2002 2022
rect 2086 2018 2090 2022
rect 2158 2018 2162 2022
rect 2198 2018 2202 2022
rect 2254 2018 2258 2022
rect 2518 2018 2522 2022
rect 3118 2018 3122 2022
rect 3238 2018 3242 2022
rect 3494 2018 3498 2022
rect 3510 2018 3514 2022
rect 482 2003 486 2007
rect 489 2003 493 2007
rect 1514 2003 1518 2007
rect 1521 2003 1525 2007
rect 2538 2003 2542 2007
rect 2545 2003 2549 2007
rect 654 1988 658 1992
rect 806 1988 810 1992
rect 1374 1988 1378 1992
rect 1406 1988 1410 1992
rect 1598 1988 1602 1992
rect 1678 1988 1682 1992
rect 1750 1988 1754 1992
rect 1870 1988 1874 1992
rect 1910 1988 1914 1992
rect 1950 1988 1954 1992
rect 2038 1988 2042 1992
rect 2166 1988 2170 1992
rect 2214 1988 2218 1992
rect 2270 1988 2274 1992
rect 2382 1988 2386 1992
rect 2422 1988 2426 1992
rect 2446 1988 2450 1992
rect 2470 1988 2474 1992
rect 2518 1988 2522 1992
rect 2566 1988 2570 1992
rect 2750 1988 2754 1992
rect 2806 1988 2810 1992
rect 2894 1988 2898 1992
rect 2942 1988 2946 1992
rect 2990 1988 2994 1992
rect 3470 1988 3474 1992
rect 70 1968 74 1972
rect 766 1968 770 1972
rect 1022 1968 1026 1972
rect 1102 1968 1106 1972
rect 1726 1968 1730 1972
rect 1734 1968 1738 1972
rect 1862 1968 1866 1972
rect 1958 1968 1962 1972
rect 2198 1968 2202 1972
rect 2262 1968 2266 1972
rect 2742 1968 2746 1972
rect 3462 1968 3466 1972
rect 3478 1968 3482 1972
rect 3518 1968 3522 1972
rect 14 1948 18 1952
rect 94 1948 98 1952
rect 206 1958 210 1962
rect 246 1958 250 1962
rect 286 1958 290 1962
rect 374 1958 378 1962
rect 382 1958 386 1962
rect 422 1958 426 1962
rect 430 1958 434 1962
rect 502 1958 506 1962
rect 534 1958 538 1962
rect 566 1958 570 1962
rect 590 1958 594 1962
rect 614 1958 618 1962
rect 670 1958 674 1962
rect 726 1958 730 1962
rect 734 1958 738 1962
rect 782 1958 786 1962
rect 822 1958 826 1962
rect 878 1958 882 1962
rect 886 1958 890 1962
rect 958 1958 962 1962
rect 966 1958 970 1962
rect 1038 1958 1042 1962
rect 1062 1958 1066 1962
rect 134 1948 138 1952
rect 166 1948 170 1952
rect 174 1948 178 1952
rect 190 1948 194 1952
rect 238 1948 242 1952
rect 270 1948 274 1952
rect 310 1948 314 1952
rect 342 1948 346 1952
rect 350 1948 354 1952
rect 478 1948 482 1952
rect 526 1948 530 1952
rect 550 1948 554 1952
rect 630 1948 634 1952
rect 654 1948 658 1952
rect 670 1948 674 1952
rect 710 1948 714 1952
rect 766 1948 770 1952
rect 790 1948 794 1952
rect 846 1948 850 1952
rect 926 1948 930 1952
rect 1022 1948 1026 1952
rect 1078 1948 1082 1952
rect 1126 1958 1130 1962
rect 1166 1958 1170 1962
rect 1182 1948 1186 1952
rect 1190 1948 1194 1952
rect 1206 1948 1210 1952
rect 1238 1958 1242 1962
rect 1286 1958 1290 1962
rect 1318 1958 1322 1962
rect 1350 1958 1354 1962
rect 1358 1958 1362 1962
rect 1390 1958 1394 1962
rect 1438 1958 1442 1962
rect 1478 1958 1482 1962
rect 1526 1958 1530 1962
rect 1686 1958 1690 1962
rect 1718 1958 1722 1962
rect 1782 1958 1786 1962
rect 1846 1958 1850 1962
rect 1878 1958 1882 1962
rect 1942 1958 1946 1962
rect 2054 1958 2058 1962
rect 2110 1958 2114 1962
rect 2142 1958 2146 1962
rect 2182 1958 2186 1962
rect 2278 1958 2282 1962
rect 2366 1958 2370 1962
rect 2398 1958 2402 1962
rect 2582 1958 2586 1962
rect 2710 1958 2714 1962
rect 2758 1958 2762 1962
rect 2846 1958 2850 1962
rect 2862 1958 2866 1962
rect 2950 1958 2954 1962
rect 3006 1958 3010 1962
rect 3126 1958 3130 1962
rect 3166 1958 3170 1962
rect 3198 1958 3202 1962
rect 3246 1958 3250 1962
rect 3262 1958 3266 1962
rect 3422 1958 3426 1962
rect 3430 1958 3434 1962
rect 1270 1948 1274 1952
rect 1302 1948 1306 1952
rect 1326 1948 1330 1952
rect 1374 1948 1378 1952
rect 1406 1948 1410 1952
rect 1470 1948 1474 1952
rect 1494 1948 1498 1952
rect 1542 1948 1546 1952
rect 1550 1948 1554 1952
rect 1598 1948 1602 1952
rect 1646 1948 1650 1952
rect 1654 1948 1658 1952
rect 1694 1948 1698 1952
rect 1702 1948 1706 1952
rect 1726 1948 1730 1952
rect 1798 1948 1802 1952
rect 1838 1948 1842 1952
rect 1854 1948 1858 1952
rect 1894 1948 1898 1952
rect 1934 1948 1938 1952
rect 1950 1948 1954 1952
rect 1990 1948 1994 1952
rect 2038 1948 2042 1952
rect 2078 1948 2082 1952
rect 2086 1948 2090 1952
rect 2166 1948 2170 1952
rect 2198 1948 2202 1952
rect 2230 1948 2234 1952
rect 2246 1948 2250 1952
rect 2270 1948 2274 1952
rect 2318 1948 2322 1952
rect 2350 1948 2354 1952
rect 2382 1948 2386 1952
rect 2406 1948 2410 1952
rect 2462 1948 2466 1952
rect 2486 1948 2490 1952
rect 2550 1948 2554 1952
rect 2566 1948 2570 1952
rect 2606 1948 2610 1952
rect 2614 1948 2618 1952
rect 2638 1948 2642 1952
rect 2646 1948 2650 1952
rect 2678 1948 2682 1952
rect 2750 1948 2754 1952
rect 2766 1948 2770 1952
rect 2814 1948 2818 1952
rect 2870 1948 2874 1952
rect 2918 1948 2922 1952
rect 2958 1948 2962 1952
rect 2966 1948 2970 1952
rect 2990 1948 2994 1952
rect 3014 1948 3018 1952
rect 3054 1948 3058 1952
rect 3086 1948 3090 1952
rect 3102 1948 3106 1952
rect 3134 1948 3138 1952
rect 3142 1948 3146 1952
rect 3182 1948 3186 1952
rect 3238 1948 3242 1952
rect 3270 1948 3274 1952
rect 3286 1948 3290 1952
rect 3302 1948 3306 1952
rect 3326 1948 3330 1952
rect 6 1938 10 1942
rect 38 1938 42 1942
rect 86 1938 90 1942
rect 102 1938 106 1942
rect 126 1938 130 1942
rect 182 1938 186 1942
rect 230 1938 234 1942
rect 270 1938 274 1942
rect 398 1938 402 1942
rect 406 1938 410 1942
rect 446 1938 450 1942
rect 478 1938 482 1942
rect 526 1938 530 1942
rect 542 1938 546 1942
rect 566 1938 570 1942
rect 582 1938 586 1942
rect 606 1938 610 1942
rect 622 1938 626 1942
rect 638 1938 642 1942
rect 694 1938 698 1942
rect 750 1938 754 1942
rect 758 1938 762 1942
rect 846 1938 850 1942
rect 854 1938 858 1942
rect 870 1938 874 1942
rect 902 1938 906 1942
rect 934 1938 938 1942
rect 942 1938 946 1942
rect 982 1938 986 1942
rect 1030 1938 1034 1942
rect 1054 1938 1058 1942
rect 1086 1938 1090 1942
rect 1094 1938 1098 1942
rect 1142 1938 1146 1942
rect 1198 1938 1202 1942
rect 1206 1938 1210 1942
rect 1254 1938 1258 1942
rect 1294 1938 1298 1942
rect 1326 1938 1330 1942
rect 1382 1938 1386 1942
rect 1414 1938 1418 1942
rect 1422 1938 1426 1942
rect 1438 1938 1442 1942
rect 1462 1938 1466 1942
rect 1502 1938 1506 1942
rect 1534 1938 1538 1942
rect 1550 1938 1554 1942
rect 1574 1938 1578 1942
rect 1590 1938 1594 1942
rect 1638 1938 1642 1942
rect 1654 1938 1658 1942
rect 1710 1938 1714 1942
rect 1766 1938 1770 1942
rect 1814 1938 1818 1942
rect 1830 1938 1834 1942
rect 1902 1938 1906 1942
rect 1926 1938 1930 1942
rect 2030 1938 2034 1942
rect 2086 1938 2090 1942
rect 2094 1938 2098 1942
rect 2126 1938 2130 1942
rect 2158 1938 2162 1942
rect 2238 1938 2242 1942
rect 2294 1938 2298 1942
rect 2342 1938 2346 1942
rect 2374 1938 2378 1942
rect 2478 1938 2482 1942
rect 2558 1938 2562 1942
rect 3358 1947 3362 1951
rect 3390 1948 3394 1952
rect 3454 1948 3458 1952
rect 3502 1948 3506 1952
rect 3526 1948 3530 1952
rect 2686 1938 2690 1942
rect 2726 1938 2730 1942
rect 2774 1938 2778 1942
rect 2822 1938 2826 1942
rect 2846 1938 2850 1942
rect 2878 1938 2882 1942
rect 2926 1938 2930 1942
rect 2974 1938 2978 1942
rect 2982 1938 2986 1942
rect 3038 1938 3042 1942
rect 3094 1938 3098 1942
rect 3150 1938 3154 1942
rect 3174 1938 3178 1942
rect 3214 1938 3218 1942
rect 3238 1938 3242 1942
rect 3270 1938 3274 1942
rect 3294 1938 3298 1942
rect 3310 1938 3314 1942
rect 3342 1938 3346 1942
rect 3478 1938 3482 1942
rect 3558 1938 3562 1942
rect 70 1928 74 1932
rect 158 1928 162 1932
rect 302 1928 306 1932
rect 694 1928 698 1932
rect 1446 1928 1450 1932
rect 1558 1928 1562 1932
rect 1622 1928 1626 1932
rect 1678 1928 1682 1932
rect 1774 1928 1778 1932
rect 1814 1928 1818 1932
rect 1910 1928 1914 1932
rect 1974 1928 1978 1932
rect 2062 1928 2066 1932
rect 2102 1928 2106 1932
rect 2134 1928 2138 1932
rect 2142 1928 2146 1932
rect 2222 1928 2226 1932
rect 2286 1928 2290 1932
rect 2334 1928 2338 1932
rect 2502 1928 2506 1932
rect 2590 1928 2594 1932
rect 2662 1928 2666 1932
rect 2702 1928 2706 1932
rect 2790 1928 2794 1932
rect 2798 1928 2802 1932
rect 2838 1928 2842 1932
rect 2910 1928 2914 1932
rect 2942 1928 2946 1932
rect 3030 1928 3034 1932
rect 3070 1928 3074 1932
rect 3110 1928 3114 1932
rect 3118 1928 3122 1932
rect 3166 1928 3170 1932
rect 3230 1928 3234 1932
rect 3310 1928 3314 1932
rect 3494 1928 3498 1932
rect 30 1918 34 1922
rect 110 1918 114 1922
rect 222 1918 226 1922
rect 246 1918 250 1922
rect 286 1918 290 1922
rect 294 1918 298 1922
rect 326 1918 330 1922
rect 366 1918 370 1922
rect 390 1918 394 1922
rect 422 1918 426 1922
rect 454 1918 458 1922
rect 502 1918 506 1922
rect 566 1918 570 1922
rect 590 1918 594 1922
rect 686 1918 690 1922
rect 726 1918 730 1922
rect 742 1918 746 1922
rect 822 1918 826 1922
rect 910 1918 914 1922
rect 950 1918 954 1922
rect 1046 1918 1050 1922
rect 1062 1918 1066 1922
rect 1230 1918 1234 1922
rect 1286 1918 1290 1922
rect 1318 1918 1322 1922
rect 1350 1918 1354 1922
rect 1438 1918 1442 1922
rect 1478 1918 1482 1922
rect 1782 1918 1786 1922
rect 1822 1918 1826 1922
rect 1878 1918 1882 1922
rect 2310 1918 2314 1922
rect 2326 1918 2330 1922
rect 2494 1918 2498 1922
rect 2598 1918 2602 1922
rect 2694 1918 2698 1922
rect 2710 1918 2714 1922
rect 2782 1918 2786 1922
rect 2862 1918 2866 1922
rect 3222 1918 3226 1922
rect 994 1903 998 1907
rect 1001 1903 1005 1907
rect 2026 1903 2030 1907
rect 2033 1903 2037 1907
rect 3042 1903 3046 1907
rect 3049 1903 3053 1907
rect 1326 1888 1330 1892
rect 1342 1888 1346 1892
rect 1414 1888 1418 1892
rect 1486 1888 1490 1892
rect 1582 1888 1586 1892
rect 1662 1888 1666 1892
rect 1718 1888 1722 1892
rect 1750 1888 1754 1892
rect 1782 1888 1786 1892
rect 1870 1888 1874 1892
rect 1934 1888 1938 1892
rect 2062 1888 2066 1892
rect 2094 1888 2098 1892
rect 2190 1888 2194 1892
rect 2214 1888 2218 1892
rect 2254 1888 2258 1892
rect 2278 1888 2282 1892
rect 2318 1888 2322 1892
rect 2454 1888 2458 1892
rect 2494 1888 2498 1892
rect 2510 1888 2514 1892
rect 2854 1888 2858 1892
rect 2886 1888 2890 1892
rect 2918 1888 2922 1892
rect 3014 1888 3018 1892
rect 3086 1888 3090 1892
rect 3118 1888 3122 1892
rect 3382 1888 3386 1892
rect 3510 1888 3514 1892
rect 3518 1888 3522 1892
rect 94 1878 98 1882
rect 102 1878 106 1882
rect 142 1878 146 1882
rect 214 1878 218 1882
rect 478 1878 482 1882
rect 510 1878 514 1882
rect 526 1878 530 1882
rect 606 1878 610 1882
rect 678 1878 682 1882
rect 902 1878 906 1882
rect 966 1878 970 1882
rect 1062 1878 1066 1882
rect 1142 1878 1146 1882
rect 1390 1878 1394 1882
rect 1422 1878 1426 1882
rect 1478 1878 1482 1882
rect 1550 1878 1554 1882
rect 1646 1878 1650 1882
rect 1942 1878 1946 1882
rect 1982 1878 1986 1882
rect 1990 1878 1994 1882
rect 2030 1878 2034 1882
rect 2038 1878 2042 1882
rect 2118 1878 2122 1882
rect 2182 1878 2186 1882
rect 2238 1878 2242 1882
rect 2246 1878 2250 1882
rect 2326 1878 2330 1882
rect 2622 1878 2626 1882
rect 2654 1878 2658 1882
rect 2662 1878 2666 1882
rect 2686 1878 2690 1882
rect 2814 1878 2818 1882
rect 2862 1878 2866 1882
rect 2878 1878 2882 1882
rect 3022 1878 3026 1882
rect 3094 1878 3098 1882
rect 3110 1878 3114 1882
rect 3230 1878 3234 1882
rect 3446 1878 3450 1882
rect 3526 1878 3530 1882
rect 6 1868 10 1872
rect 150 1868 154 1872
rect 294 1868 298 1872
rect 342 1868 346 1872
rect 350 1868 354 1872
rect 422 1868 426 1872
rect 534 1868 538 1872
rect 590 1868 594 1872
rect 614 1868 618 1872
rect 662 1868 666 1872
rect 710 1868 714 1872
rect 742 1868 746 1872
rect 766 1868 770 1872
rect 838 1868 842 1872
rect 870 1868 874 1872
rect 942 1868 946 1872
rect 998 1868 1002 1872
rect 1014 1868 1018 1872
rect 1086 1868 1090 1872
rect 1118 1868 1122 1872
rect 1214 1868 1218 1872
rect 1318 1868 1322 1872
rect 1358 1868 1362 1872
rect 1374 1868 1378 1872
rect 1494 1868 1498 1872
rect 1518 1868 1522 1872
rect 1590 1868 1594 1872
rect 1630 1868 1634 1872
rect 1638 1868 1642 1872
rect 1670 1868 1674 1872
rect 1678 1868 1682 1872
rect 1710 1868 1714 1872
rect 1750 1868 1754 1872
rect 1766 1868 1770 1872
rect 1774 1868 1778 1872
rect 1830 1868 1834 1872
rect 1846 1868 1850 1872
rect 1862 1868 1866 1872
rect 1886 1868 1890 1872
rect 1894 1868 1898 1872
rect 1950 1868 1954 1872
rect 1982 1868 1986 1872
rect 1998 1868 2002 1872
rect 2046 1868 2050 1872
rect 2086 1868 2090 1872
rect 2118 1868 2122 1872
rect 2134 1868 2138 1872
rect 2150 1868 2154 1872
rect 2166 1868 2170 1872
rect 2198 1868 2202 1872
rect 2230 1868 2234 1872
rect 2262 1868 2266 1872
rect 2294 1868 2298 1872
rect 2310 1868 2314 1872
rect 2334 1868 2338 1872
rect 2350 1868 2354 1872
rect 2358 1868 2362 1872
rect 2390 1868 2394 1872
rect 2430 1868 2434 1872
rect 2446 1868 2450 1872
rect 2486 1868 2490 1872
rect 2526 1868 2530 1872
rect 2646 1868 2650 1872
rect 2662 1868 2666 1872
rect 2678 1868 2682 1872
rect 2710 1868 2714 1872
rect 2750 1868 2754 1872
rect 2790 1868 2794 1872
rect 2846 1868 2850 1872
rect 2862 1868 2866 1872
rect 2918 1868 2922 1872
rect 2934 1868 2938 1872
rect 2942 1868 2946 1872
rect 2990 1868 2994 1872
rect 3006 1868 3010 1872
rect 3078 1868 3082 1872
rect 3142 1868 3146 1872
rect 3150 1868 3154 1872
rect 3174 1868 3178 1872
rect 3222 1868 3226 1872
rect 3246 1868 3250 1872
rect 3270 1868 3274 1872
rect 3286 1868 3290 1872
rect 3390 1868 3394 1872
rect 30 1858 34 1862
rect 46 1858 50 1862
rect 70 1858 74 1862
rect 78 1858 82 1862
rect 118 1858 122 1862
rect 182 1858 186 1862
rect 190 1858 194 1862
rect 222 1858 226 1862
rect 230 1858 234 1862
rect 254 1858 258 1862
rect 294 1858 298 1862
rect 310 1858 314 1862
rect 334 1858 338 1862
rect 374 1858 378 1862
rect 382 1858 386 1862
rect 430 1858 434 1862
rect 454 1858 458 1862
rect 462 1858 466 1862
rect 534 1858 538 1862
rect 550 1858 554 1862
rect 582 1858 586 1862
rect 654 1858 658 1862
rect 782 1858 786 1862
rect 798 1858 802 1862
rect 822 1858 826 1862
rect 846 1858 850 1862
rect 862 1858 866 1862
rect 918 1858 922 1862
rect 926 1858 930 1862
rect 1030 1858 1034 1862
rect 1038 1858 1042 1862
rect 1102 1858 1106 1862
rect 1110 1858 1114 1862
rect 1126 1858 1130 1862
rect 1134 1858 1138 1862
rect 1158 1858 1162 1862
rect 1174 1858 1178 1862
rect 1182 1858 1186 1862
rect 1206 1858 1210 1862
rect 1222 1858 1226 1862
rect 1254 1858 1258 1862
rect 1262 1858 1266 1862
rect 1278 1858 1282 1862
rect 1302 1858 1306 1862
rect 1366 1858 1370 1862
rect 1398 1858 1402 1862
rect 1430 1858 1434 1862
rect 1438 1858 1442 1862
rect 1462 1858 1466 1862
rect 1502 1858 1506 1862
rect 1526 1858 1530 1862
rect 1566 1858 1570 1862
rect 1598 1858 1602 1862
rect 1614 1858 1618 1862
rect 1622 1858 1626 1862
rect 1678 1858 1682 1862
rect 1702 1858 1706 1862
rect 1718 1858 1722 1862
rect 1734 1858 1738 1862
rect 1798 1858 1802 1862
rect 1822 1858 1826 1862
rect 1838 1858 1842 1862
rect 1862 1858 1866 1862
rect 1918 1858 1922 1862
rect 1958 1858 1962 1862
rect 2006 1858 2010 1862
rect 2014 1858 2018 1862
rect 2078 1858 2082 1862
rect 2110 1858 2114 1862
rect 2142 1858 2146 1862
rect 2158 1858 2162 1862
rect 2206 1858 2210 1862
rect 2270 1858 2274 1862
rect 2302 1858 2306 1862
rect 2574 1858 2578 1862
rect 2606 1858 2610 1862
rect 2622 1858 2626 1862
rect 2638 1858 2642 1862
rect 2678 1858 2682 1862
rect 2702 1858 2706 1862
rect 2710 1858 2714 1862
rect 2742 1858 2746 1862
rect 2758 1858 2762 1862
rect 2830 1858 2834 1862
rect 2838 1858 2842 1862
rect 2902 1858 2906 1862
rect 2998 1858 3002 1862
rect 3070 1858 3074 1862
rect 3110 1858 3114 1862
rect 3142 1858 3146 1862
rect 3238 1858 3242 1862
rect 3254 1858 3258 1862
rect 3278 1858 3282 1862
rect 3318 1859 3322 1863
rect 3342 1858 3346 1862
rect 3398 1858 3402 1862
rect 3414 1858 3418 1862
rect 3446 1859 3450 1863
rect 3526 1858 3530 1862
rect 102 1848 106 1852
rect 166 1848 170 1852
rect 246 1848 250 1852
rect 270 1848 274 1852
rect 366 1848 370 1852
rect 558 1848 562 1852
rect 566 1848 570 1852
rect 630 1848 634 1852
rect 686 1848 690 1852
rect 718 1848 722 1852
rect 742 1848 746 1852
rect 758 1848 762 1852
rect 782 1848 786 1852
rect 958 1848 962 1852
rect 982 1848 986 1852
rect 1046 1848 1050 1852
rect 1334 1848 1338 1852
rect 1342 1848 1346 1852
rect 1582 1848 1586 1852
rect 1654 1848 1658 1852
rect 1702 1848 1706 1852
rect 1750 1848 1754 1852
rect 1790 1848 1794 1852
rect 1822 1848 1826 1852
rect 1870 1848 1874 1852
rect 1910 1848 1914 1852
rect 1974 1848 1978 1852
rect 2174 1848 2178 1852
rect 2278 1848 2282 1852
rect 2582 1848 2586 1852
rect 2590 1848 2594 1852
rect 2734 1848 2738 1852
rect 2774 1848 2778 1852
rect 2918 1848 2922 1852
rect 3030 1848 3034 1852
rect 3118 1848 3122 1852
rect 3166 1848 3170 1852
rect 3206 1848 3210 1852
rect 3262 1848 3266 1852
rect 3414 1848 3418 1852
rect 734 1838 738 1842
rect 1070 1838 1074 1842
rect 1286 1838 1290 1842
rect 2566 1838 2570 1842
rect 2606 1838 2610 1842
rect 2702 1838 2706 1842
rect 2958 1838 2962 1842
rect 3558 1838 3562 1842
rect 518 1828 522 1832
rect 62 1818 66 1822
rect 86 1818 90 1822
rect 358 1818 362 1822
rect 438 1818 442 1822
rect 470 1818 474 1822
rect 502 1818 506 1822
rect 582 1818 586 1822
rect 598 1818 602 1822
rect 654 1818 658 1822
rect 670 1818 674 1822
rect 702 1818 706 1822
rect 774 1818 778 1822
rect 814 1818 818 1822
rect 974 1818 978 1822
rect 990 1818 994 1822
rect 1190 1818 1194 1822
rect 1446 1818 1450 1822
rect 2414 1818 2418 1822
rect 2438 1818 2442 1822
rect 2494 1818 2498 1822
rect 2598 1818 2602 1822
rect 2718 1818 2722 1822
rect 2798 1818 2802 1822
rect 3158 1818 3162 1822
rect 482 1803 486 1807
rect 489 1803 493 1807
rect 1514 1803 1518 1807
rect 1521 1803 1525 1807
rect 2538 1803 2542 1807
rect 2545 1803 2549 1807
rect 190 1788 194 1792
rect 590 1788 594 1792
rect 1174 1788 1178 1792
rect 1198 1788 1202 1792
rect 1446 1788 1450 1792
rect 1486 1788 1490 1792
rect 1598 1788 1602 1792
rect 1662 1788 1666 1792
rect 1782 1788 1786 1792
rect 1854 1788 1858 1792
rect 2054 1788 2058 1792
rect 2110 1788 2114 1792
rect 2158 1788 2162 1792
rect 2254 1788 2258 1792
rect 2310 1788 2314 1792
rect 2654 1788 2658 1792
rect 2678 1788 2682 1792
rect 2758 1788 2762 1792
rect 2790 1788 2794 1792
rect 2990 1788 2994 1792
rect 3150 1788 3154 1792
rect 3278 1788 3282 1792
rect 3366 1788 3370 1792
rect 3398 1788 3402 1792
rect 718 1778 722 1782
rect 1134 1778 1138 1782
rect 1390 1778 1394 1782
rect 1726 1778 1730 1782
rect 1822 1778 1826 1782
rect 1926 1778 1930 1782
rect 2334 1778 2338 1782
rect 3230 1778 3234 1782
rect 1286 1768 1290 1772
rect 1454 1768 1458 1772
rect 2494 1768 2498 1772
rect 2718 1768 2722 1772
rect 6 1758 10 1762
rect 38 1758 42 1762
rect 62 1758 66 1762
rect 110 1758 114 1762
rect 134 1758 138 1762
rect 142 1758 146 1762
rect 206 1758 210 1762
rect 254 1758 258 1762
rect 286 1758 290 1762
rect 310 1758 314 1762
rect 358 1758 362 1762
rect 382 1758 386 1762
rect 414 1758 418 1762
rect 526 1758 530 1762
rect 622 1758 626 1762
rect 630 1758 634 1762
rect 22 1748 26 1752
rect 78 1748 82 1752
rect 94 1748 98 1752
rect 158 1748 162 1752
rect 174 1748 178 1752
rect 198 1748 202 1752
rect 222 1748 226 1752
rect 270 1748 274 1752
rect 350 1748 354 1752
rect 398 1748 402 1752
rect 430 1748 434 1752
rect 446 1748 450 1752
rect 454 1748 458 1752
rect 478 1748 482 1752
rect 534 1748 538 1752
rect 566 1748 570 1752
rect 606 1748 610 1752
rect 646 1748 650 1752
rect 662 1748 666 1752
rect 686 1758 690 1762
rect 734 1758 738 1762
rect 798 1758 802 1762
rect 806 1758 810 1762
rect 822 1758 826 1762
rect 910 1758 914 1762
rect 918 1758 922 1762
rect 958 1758 962 1762
rect 982 1758 986 1762
rect 1030 1758 1034 1762
rect 1054 1758 1058 1762
rect 710 1748 714 1752
rect 742 1748 746 1752
rect 766 1748 770 1752
rect 878 1748 882 1752
rect 1014 1748 1018 1752
rect 1094 1758 1098 1762
rect 1166 1758 1170 1762
rect 1302 1758 1306 1762
rect 1358 1758 1362 1762
rect 1438 1758 1442 1762
rect 1470 1758 1474 1762
rect 1518 1758 1522 1762
rect 1534 1758 1538 1762
rect 1550 1758 1554 1762
rect 1582 1758 1586 1762
rect 1614 1758 1618 1762
rect 1654 1758 1658 1762
rect 1702 1758 1706 1762
rect 1710 1758 1714 1762
rect 1766 1758 1770 1762
rect 1910 1758 1914 1762
rect 2126 1758 2130 1762
rect 2190 1758 2194 1762
rect 2270 1758 2274 1762
rect 2302 1758 2306 1762
rect 2662 1758 2666 1762
rect 2718 1758 2722 1762
rect 2894 1758 2898 1762
rect 3094 1758 3098 1762
rect 3166 1758 3170 1762
rect 3206 1758 3210 1762
rect 3254 1758 3258 1762
rect 3294 1758 3298 1762
rect 3358 1758 3362 1762
rect 3382 1758 3386 1762
rect 3510 1758 3514 1762
rect 1078 1748 1082 1752
rect 1150 1748 1154 1752
rect 1190 1748 1194 1752
rect 1214 1748 1218 1752
rect 1222 1748 1226 1752
rect 1246 1748 1250 1752
rect 1262 1748 1266 1752
rect 1278 1748 1282 1752
rect 1310 1748 1314 1752
rect 1350 1748 1354 1752
rect 1366 1748 1370 1752
rect 1374 1748 1378 1752
rect 1398 1748 1402 1752
rect 1422 1748 1426 1752
rect 1462 1748 1466 1752
rect 1486 1748 1490 1752
rect 1510 1748 1514 1752
rect 1566 1748 1570 1752
rect 1582 1748 1586 1752
rect 1598 1748 1602 1752
rect 1622 1748 1626 1752
rect 1638 1748 1642 1752
rect 1678 1748 1682 1752
rect 1726 1748 1730 1752
rect 1742 1748 1746 1752
rect 1798 1748 1802 1752
rect 1830 1748 1834 1752
rect 1846 1748 1850 1752
rect 1862 1748 1866 1752
rect 1870 1748 1874 1752
rect 1902 1748 1906 1752
rect 1926 1748 1930 1752
rect 1982 1748 1986 1752
rect 1998 1748 2002 1752
rect 2046 1748 2050 1752
rect 2062 1748 2066 1752
rect 2078 1748 2082 1752
rect 2102 1748 2106 1752
rect 2126 1748 2130 1752
rect 2150 1748 2154 1752
rect 2174 1748 2178 1752
rect 2222 1748 2226 1752
rect 2254 1748 2258 1752
rect 2286 1748 2290 1752
rect 2350 1748 2354 1752
rect 2366 1748 2370 1752
rect 2414 1748 2418 1752
rect 2446 1748 2450 1752
rect 2542 1748 2546 1752
rect 2574 1748 2578 1752
rect 2654 1748 2658 1752
rect 2678 1748 2682 1752
rect 2790 1748 2794 1752
rect 2814 1748 2818 1752
rect 2878 1748 2882 1752
rect 2902 1748 2906 1752
rect 2934 1748 2938 1752
rect 2958 1748 2962 1752
rect 3030 1748 3034 1752
rect 3070 1748 3074 1752
rect 3110 1748 3114 1752
rect 3150 1748 3154 1752
rect 3262 1748 3266 1752
rect 3350 1748 3354 1752
rect 3398 1748 3402 1752
rect 3494 1748 3498 1752
rect 3542 1748 3546 1752
rect 30 1738 34 1742
rect 38 1738 42 1742
rect 54 1738 58 1742
rect 86 1738 90 1742
rect 118 1738 122 1742
rect 150 1738 154 1742
rect 166 1738 170 1742
rect 230 1738 234 1742
rect 238 1738 242 1742
rect 262 1738 266 1742
rect 294 1738 298 1742
rect 374 1738 378 1742
rect 406 1738 410 1742
rect 422 1738 426 1742
rect 438 1738 442 1742
rect 494 1738 498 1742
rect 510 1738 514 1742
rect 542 1738 546 1742
rect 590 1738 594 1742
rect 606 1738 610 1742
rect 646 1738 650 1742
rect 702 1738 706 1742
rect 710 1738 714 1742
rect 774 1738 778 1742
rect 822 1738 826 1742
rect 846 1738 850 1742
rect 878 1738 882 1742
rect 886 1738 890 1742
rect 934 1738 938 1742
rect 942 1738 946 1742
rect 958 1738 962 1742
rect 966 1738 970 1742
rect 982 1738 986 1742
rect 1038 1738 1042 1742
rect 1086 1738 1090 1742
rect 1110 1738 1114 1742
rect 1142 1738 1146 1742
rect 1150 1738 1154 1742
rect 1286 1738 1290 1742
rect 1334 1738 1338 1742
rect 1414 1738 1418 1742
rect 1430 1738 1434 1742
rect 1478 1738 1482 1742
rect 1526 1738 1530 1742
rect 1558 1738 1562 1742
rect 1590 1738 1594 1742
rect 1630 1738 1634 1742
rect 1670 1738 1674 1742
rect 1678 1738 1682 1742
rect 1742 1738 1746 1742
rect 1774 1738 1778 1742
rect 1814 1738 1818 1742
rect 1838 1738 1842 1742
rect 1894 1738 1898 1742
rect 1958 1738 1962 1742
rect 1990 1738 1994 1742
rect 2038 1738 2042 1742
rect 2070 1738 2074 1742
rect 2086 1738 2090 1742
rect 2150 1738 2154 1742
rect 2166 1738 2170 1742
rect 2198 1738 2202 1742
rect 2214 1738 2218 1742
rect 2278 1738 2282 1742
rect 2358 1738 2362 1742
rect 2406 1738 2410 1742
rect 2470 1738 2474 1742
rect 2598 1738 2602 1742
rect 2686 1738 2690 1742
rect 2734 1738 2738 1742
rect 2878 1738 2882 1742
rect 2974 1738 2978 1742
rect 2998 1738 3002 1742
rect 3062 1738 3066 1742
rect 3142 1738 3146 1742
rect 3182 1738 3186 1742
rect 3206 1738 3210 1742
rect 3222 1738 3226 1742
rect 3270 1738 3274 1742
rect 3302 1738 3306 1742
rect 3350 1738 3354 1742
rect 3374 1738 3378 1742
rect 3406 1738 3410 1742
rect 3414 1738 3418 1742
rect 3486 1738 3490 1742
rect 3534 1738 3538 1742
rect 3558 1738 3562 1742
rect 318 1728 322 1732
rect 334 1728 338 1732
rect 558 1728 562 1732
rect 1062 1728 1066 1732
rect 1182 1728 1186 1732
rect 1206 1728 1210 1732
rect 1230 1728 1234 1732
rect 1278 1728 1282 1732
rect 1326 1728 1330 1732
rect 1646 1728 1650 1732
rect 1814 1728 1818 1732
rect 1878 1728 1882 1732
rect 1942 1728 1946 1732
rect 2102 1728 2106 1732
rect 2118 1728 2122 1732
rect 2150 1728 2154 1732
rect 2230 1728 2234 1732
rect 2302 1728 2306 1732
rect 2318 1728 2322 1732
rect 2390 1728 2394 1732
rect 2454 1728 2458 1732
rect 2510 1728 2514 1732
rect 2566 1728 2570 1732
rect 2590 1728 2594 1732
rect 2638 1728 2642 1732
rect 2694 1728 2698 1732
rect 2750 1728 2754 1732
rect 2782 1728 2786 1732
rect 2806 1728 2810 1732
rect 2830 1728 2834 1732
rect 2838 1728 2842 1732
rect 2854 1728 2858 1732
rect 2942 1728 2946 1732
rect 2966 1728 2970 1732
rect 3086 1728 3090 1732
rect 3126 1728 3130 1732
rect 3198 1728 3202 1732
rect 3238 1728 3242 1732
rect 3470 1728 3474 1732
rect 3518 1728 3522 1732
rect 6 1718 10 1722
rect 62 1718 66 1722
rect 110 1718 114 1722
rect 126 1718 130 1722
rect 254 1718 258 1722
rect 286 1718 290 1722
rect 310 1718 314 1722
rect 358 1718 362 1722
rect 382 1718 386 1722
rect 518 1718 522 1722
rect 614 1718 618 1722
rect 630 1718 634 1722
rect 678 1718 682 1722
rect 798 1718 802 1722
rect 806 1718 810 1722
rect 854 1718 858 1722
rect 910 1718 914 1722
rect 918 1718 922 1722
rect 982 1718 986 1722
rect 1030 1718 1034 1722
rect 1166 1718 1170 1722
rect 1702 1718 1706 1722
rect 1950 1718 1954 1722
rect 2030 1718 2034 1722
rect 2382 1718 2386 1722
rect 2398 1718 2402 1722
rect 2430 1718 2434 1722
rect 2462 1718 2466 1722
rect 2558 1718 2562 1722
rect 2582 1718 2586 1722
rect 2606 1718 2610 1722
rect 2742 1718 2746 1722
rect 2774 1718 2778 1722
rect 2798 1718 2802 1722
rect 2822 1718 2826 1722
rect 2918 1718 2922 1722
rect 3078 1718 3082 1722
rect 3094 1718 3098 1722
rect 3190 1718 3194 1722
rect 3510 1718 3514 1722
rect 3526 1718 3530 1722
rect 3550 1718 3554 1722
rect 994 1703 998 1707
rect 1001 1703 1005 1707
rect 2026 1703 2030 1707
rect 2033 1703 2037 1707
rect 3042 1703 3046 1707
rect 3049 1703 3053 1707
rect 30 1688 34 1692
rect 126 1688 130 1692
rect 246 1688 250 1692
rect 894 1688 898 1692
rect 926 1688 930 1692
rect 1294 1688 1298 1692
rect 1382 1688 1386 1692
rect 1438 1688 1442 1692
rect 1462 1688 1466 1692
rect 1518 1688 1522 1692
rect 1574 1688 1578 1692
rect 1606 1688 1610 1692
rect 1710 1688 1714 1692
rect 1742 1688 1746 1692
rect 1830 1688 1834 1692
rect 1870 1688 1874 1692
rect 1958 1688 1962 1692
rect 2062 1688 2066 1692
rect 2094 1688 2098 1692
rect 2134 1688 2138 1692
rect 2158 1688 2162 1692
rect 2198 1688 2202 1692
rect 2230 1688 2234 1692
rect 2286 1688 2290 1692
rect 2318 1688 2322 1692
rect 2342 1688 2346 1692
rect 2374 1688 2378 1692
rect 2438 1688 2442 1692
rect 2574 1688 2578 1692
rect 2614 1688 2618 1692
rect 2670 1688 2674 1692
rect 2710 1688 2714 1692
rect 2910 1688 2914 1692
rect 3014 1688 3018 1692
rect 3166 1688 3170 1692
rect 3438 1688 3442 1692
rect 3510 1688 3514 1692
rect 598 1678 602 1682
rect 86 1668 90 1672
rect 166 1668 170 1672
rect 214 1668 218 1672
rect 294 1668 298 1672
rect 302 1668 306 1672
rect 494 1668 498 1672
rect 526 1668 530 1672
rect 550 1668 554 1672
rect 654 1678 658 1682
rect 662 1678 666 1682
rect 678 1678 682 1682
rect 886 1678 890 1682
rect 1110 1678 1114 1682
rect 1118 1678 1122 1682
rect 1134 1678 1138 1682
rect 1390 1678 1394 1682
rect 1414 1678 1418 1682
rect 1422 1678 1426 1682
rect 1446 1678 1450 1682
rect 1526 1678 1530 1682
rect 1582 1678 1586 1682
rect 1614 1678 1618 1682
rect 1662 1678 1666 1682
rect 1734 1678 1738 1682
rect 1782 1678 1786 1682
rect 1838 1678 1842 1682
rect 1966 1678 1970 1682
rect 2014 1678 2018 1682
rect 2054 1678 2058 1682
rect 2086 1678 2090 1682
rect 2142 1678 2146 1682
rect 2206 1678 2210 1682
rect 2238 1678 2242 1682
rect 2278 1678 2282 1682
rect 2334 1678 2338 1682
rect 2582 1678 2586 1682
rect 2598 1678 2602 1682
rect 2966 1678 2970 1682
rect 3006 1678 3010 1682
rect 3038 1678 3042 1682
rect 3062 1678 3066 1682
rect 3102 1678 3106 1682
rect 3110 1678 3114 1682
rect 3150 1678 3154 1682
rect 3174 1678 3178 1682
rect 3214 1678 3218 1682
rect 3318 1678 3322 1682
rect 3326 1678 3330 1682
rect 622 1668 626 1672
rect 630 1668 634 1672
rect 646 1668 650 1672
rect 686 1668 690 1672
rect 742 1668 746 1672
rect 750 1668 754 1672
rect 798 1668 802 1672
rect 806 1668 810 1672
rect 854 1668 858 1672
rect 878 1668 882 1672
rect 902 1668 906 1672
rect 934 1668 938 1672
rect 958 1668 962 1672
rect 1078 1668 1082 1672
rect 1142 1668 1146 1672
rect 1270 1668 1274 1672
rect 1326 1668 1330 1672
rect 1342 1668 1346 1672
rect 1358 1668 1362 1672
rect 1374 1668 1378 1672
rect 1406 1668 1410 1672
rect 1470 1668 1474 1672
rect 1478 1668 1482 1672
rect 1542 1668 1546 1672
rect 1566 1668 1570 1672
rect 1598 1668 1602 1672
rect 1662 1668 1666 1672
rect 1686 1668 1690 1672
rect 1702 1668 1706 1672
rect 1726 1668 1730 1672
rect 1758 1668 1762 1672
rect 1822 1668 1826 1672
rect 1846 1668 1850 1672
rect 1878 1668 1882 1672
rect 1886 1668 1890 1672
rect 1918 1668 1922 1672
rect 1934 1668 1938 1672
rect 1950 1668 1954 1672
rect 1966 1668 1970 1672
rect 1990 1668 1994 1672
rect 2078 1668 2082 1672
rect 2102 1668 2106 1672
rect 2126 1668 2130 1672
rect 2166 1668 2170 1672
rect 2190 1668 2194 1672
rect 2222 1668 2226 1672
rect 2246 1668 2250 1672
rect 2262 1668 2266 1672
rect 2294 1668 2298 1672
rect 2310 1668 2314 1672
rect 2350 1668 2354 1672
rect 2366 1668 2370 1672
rect 2398 1668 2402 1672
rect 2430 1668 2434 1672
rect 2454 1668 2458 1672
rect 2462 1668 2466 1672
rect 2494 1668 2498 1672
rect 2502 1668 2506 1672
rect 2550 1668 2554 1672
rect 3446 1678 3450 1682
rect 3454 1678 3458 1682
rect 3502 1678 3506 1682
rect 3534 1678 3538 1682
rect 2622 1668 2626 1672
rect 2678 1668 2682 1672
rect 2686 1668 2690 1672
rect 2718 1668 2722 1672
rect 2750 1668 2754 1672
rect 2942 1668 2946 1672
rect 2950 1668 2954 1672
rect 2982 1668 2986 1672
rect 3198 1668 3202 1672
rect 3262 1668 3266 1672
rect 3278 1668 3282 1672
rect 3302 1668 3306 1672
rect 3342 1668 3346 1672
rect 3358 1668 3362 1672
rect 3366 1668 3370 1672
rect 3382 1668 3386 1672
rect 3414 1668 3418 1672
rect 3430 1668 3434 1672
rect 3454 1668 3458 1672
rect 3478 1668 3482 1672
rect 6 1658 10 1662
rect 38 1658 42 1662
rect 46 1658 50 1662
rect 70 1658 74 1662
rect 110 1658 114 1662
rect 206 1658 210 1662
rect 222 1658 226 1662
rect 230 1658 234 1662
rect 254 1658 258 1662
rect 294 1658 298 1662
rect 310 1658 314 1662
rect 334 1658 338 1662
rect 342 1658 346 1662
rect 366 1658 370 1662
rect 374 1658 378 1662
rect 382 1658 386 1662
rect 390 1658 394 1662
rect 414 1658 418 1662
rect 430 1658 434 1662
rect 438 1658 442 1662
rect 494 1658 498 1662
rect 502 1658 506 1662
rect 558 1658 562 1662
rect 566 1658 570 1662
rect 582 1658 586 1662
rect 598 1658 602 1662
rect 622 1658 626 1662
rect 694 1658 698 1662
rect 734 1658 738 1662
rect 758 1658 762 1662
rect 838 1658 842 1662
rect 846 1658 850 1662
rect 902 1658 906 1662
rect 966 1658 970 1662
rect 974 1658 978 1662
rect 1014 1658 1018 1662
rect 1038 1658 1042 1662
rect 1054 1658 1058 1662
rect 1078 1658 1082 1662
rect 1102 1658 1106 1662
rect 1134 1658 1138 1662
rect 1174 1658 1178 1662
rect 1206 1658 1210 1662
rect 1214 1658 1218 1662
rect 1222 1658 1226 1662
rect 1230 1658 1234 1662
rect 1254 1658 1258 1662
rect 1278 1658 1282 1662
rect 1318 1658 1322 1662
rect 1350 1658 1354 1662
rect 1366 1658 1370 1662
rect 1398 1658 1402 1662
rect 1430 1658 1434 1662
rect 1486 1658 1490 1662
rect 1534 1658 1538 1662
rect 1550 1658 1554 1662
rect 1558 1658 1562 1662
rect 1590 1658 1594 1662
rect 1638 1658 1642 1662
rect 1678 1658 1682 1662
rect 1694 1658 1698 1662
rect 1758 1658 1762 1662
rect 1766 1658 1770 1662
rect 1774 1658 1778 1662
rect 1798 1658 1802 1662
rect 1814 1658 1818 1662
rect 1854 1658 1858 1662
rect 1870 1658 1874 1662
rect 1894 1658 1898 1662
rect 1918 1658 1922 1662
rect 1942 1658 1946 1662
rect 1982 1658 1986 1662
rect 1998 1658 2002 1662
rect 2038 1658 2042 1662
rect 2078 1658 2082 1662
rect 2110 1658 2114 1662
rect 2118 1658 2122 1662
rect 2174 1658 2178 1662
rect 2182 1658 2186 1662
rect 2214 1658 2218 1662
rect 2254 1658 2258 1662
rect 2302 1658 2306 1662
rect 2358 1658 2362 1662
rect 2374 1658 2378 1662
rect 2422 1658 2426 1662
rect 2470 1658 2474 1662
rect 2486 1658 2490 1662
rect 2510 1658 2514 1662
rect 2526 1658 2530 1662
rect 2558 1658 2562 1662
rect 2582 1658 2586 1662
rect 2654 1658 2658 1662
rect 2694 1658 2698 1662
rect 2726 1658 2730 1662
rect 2774 1658 2778 1662
rect 2782 1658 2786 1662
rect 2806 1658 2810 1662
rect 2838 1658 2842 1662
rect 2878 1658 2882 1662
rect 2926 1658 2930 1662
rect 2934 1658 2938 1662
rect 2958 1658 2962 1662
rect 3078 1658 3082 1662
rect 3086 1658 3090 1662
rect 3134 1658 3138 1662
rect 3150 1658 3154 1662
rect 3214 1658 3218 1662
rect 3246 1658 3250 1662
rect 3254 1658 3258 1662
rect 3294 1658 3298 1662
rect 3342 1658 3346 1662
rect 3414 1658 3418 1662
rect 3422 1658 3426 1662
rect 3470 1658 3474 1662
rect 3486 1658 3490 1662
rect 54 1648 58 1652
rect 102 1648 106 1652
rect 158 1648 162 1652
rect 182 1648 186 1652
rect 270 1648 274 1652
rect 326 1648 330 1652
rect 454 1648 458 1652
rect 502 1648 506 1652
rect 518 1648 522 1652
rect 574 1648 578 1652
rect 710 1648 714 1652
rect 718 1648 722 1652
rect 782 1648 786 1652
rect 822 1648 826 1652
rect 926 1648 930 1652
rect 934 1648 938 1652
rect 982 1648 986 1652
rect 1054 1648 1058 1652
rect 1166 1648 1170 1652
rect 1294 1648 1298 1652
rect 1318 1648 1322 1652
rect 1334 1648 1338 1652
rect 1454 1648 1458 1652
rect 1518 1648 1522 1652
rect 1622 1648 1626 1652
rect 1638 1648 1642 1652
rect 1710 1648 1714 1652
rect 1910 1648 1914 1652
rect 2270 1648 2274 1652
rect 2326 1648 2330 1652
rect 2406 1648 2410 1652
rect 2438 1648 2442 1652
rect 2542 1648 2546 1652
rect 2574 1648 2578 1652
rect 2606 1648 2610 1652
rect 2638 1648 2642 1652
rect 2662 1648 2666 1652
rect 2742 1648 2746 1652
rect 2894 1648 2898 1652
rect 2910 1648 2914 1652
rect 3046 1648 3050 1652
rect 3182 1648 3186 1652
rect 3326 1648 3330 1652
rect 3366 1648 3370 1652
rect 3390 1648 3394 1652
rect 3406 1648 3410 1652
rect 3502 1648 3506 1652
rect 3510 1648 3514 1652
rect 86 1638 90 1642
rect 206 1638 210 1642
rect 526 1638 530 1642
rect 734 1638 738 1642
rect 878 1638 882 1642
rect 358 1628 362 1632
rect 70 1618 74 1622
rect 150 1618 154 1622
rect 286 1618 290 1622
rect 406 1618 410 1622
rect 606 1618 610 1622
rect 670 1618 674 1622
rect 694 1618 698 1622
rect 758 1618 762 1622
rect 1030 1618 1034 1622
rect 1070 1618 1074 1622
rect 1086 1618 1090 1622
rect 1126 1618 1130 1622
rect 1150 1618 1154 1622
rect 1190 1618 1194 1622
rect 1246 1618 1250 1622
rect 1926 1618 1930 1622
rect 2486 1618 2490 1622
rect 2726 1618 2730 1622
rect 2822 1618 2826 1622
rect 2862 1618 2866 1622
rect 2998 1618 3002 1622
rect 3070 1618 3074 1622
rect 3086 1618 3090 1622
rect 3126 1618 3130 1622
rect 3134 1618 3138 1622
rect 3190 1618 3194 1622
rect 3230 1618 3234 1622
rect 3278 1618 3282 1622
rect 482 1603 486 1607
rect 489 1603 493 1607
rect 1514 1603 1518 1607
rect 1521 1603 1525 1607
rect 2538 1603 2542 1607
rect 2545 1603 2549 1607
rect 1238 1588 1242 1592
rect 1406 1588 1410 1592
rect 1430 1588 1434 1592
rect 1598 1588 1602 1592
rect 1670 1588 1674 1592
rect 1958 1588 1962 1592
rect 2070 1588 2074 1592
rect 2214 1588 2218 1592
rect 2238 1588 2242 1592
rect 2254 1588 2258 1592
rect 2302 1588 2306 1592
rect 2438 1588 2442 1592
rect 2486 1588 2490 1592
rect 2750 1588 2754 1592
rect 2774 1588 2778 1592
rect 2854 1588 2858 1592
rect 2990 1588 2994 1592
rect 3150 1588 3154 1592
rect 3190 1588 3194 1592
rect 3374 1588 3378 1592
rect 3502 1588 3506 1592
rect 222 1578 226 1582
rect 718 1578 722 1582
rect 878 1578 882 1582
rect 2150 1578 2154 1582
rect 3510 1578 3514 1582
rect 302 1568 306 1572
rect 414 1568 418 1572
rect 926 1568 930 1572
rect 1318 1568 1322 1572
rect 1886 1568 1890 1572
rect 2014 1568 2018 1572
rect 2478 1568 2482 1572
rect 2494 1568 2498 1572
rect 2550 1568 2554 1572
rect 2742 1568 2746 1572
rect 2806 1568 2810 1572
rect 2998 1568 3002 1572
rect 3158 1568 3162 1572
rect 3558 1568 3562 1572
rect 14 1558 18 1562
rect 54 1558 58 1562
rect 78 1558 82 1562
rect 86 1558 90 1562
rect 142 1558 146 1562
rect 150 1558 154 1562
rect 190 1558 194 1562
rect 270 1558 274 1562
rect 318 1558 322 1562
rect 398 1558 402 1562
rect 446 1558 450 1562
rect 470 1558 474 1562
rect 30 1548 34 1552
rect 102 1548 106 1552
rect 126 1548 130 1552
rect 142 1548 146 1552
rect 198 1548 202 1552
rect 206 1548 210 1552
rect 230 1548 234 1552
rect 238 1548 242 1552
rect 302 1548 306 1552
rect 318 1548 322 1552
rect 334 1548 338 1552
rect 358 1548 362 1552
rect 390 1548 394 1552
rect 414 1548 418 1552
rect 502 1548 506 1552
rect 526 1558 530 1562
rect 598 1558 602 1562
rect 630 1558 634 1562
rect 542 1548 546 1552
rect 566 1548 570 1552
rect 582 1548 586 1552
rect 614 1548 618 1552
rect 622 1548 626 1552
rect 774 1558 778 1562
rect 654 1548 658 1552
rect 662 1548 666 1552
rect 694 1548 698 1552
rect 726 1548 730 1552
rect 750 1548 754 1552
rect 830 1558 834 1562
rect 886 1558 890 1562
rect 910 1558 914 1562
rect 950 1558 954 1562
rect 982 1558 986 1562
rect 1054 1558 1058 1562
rect 1094 1558 1098 1562
rect 1134 1558 1138 1562
rect 790 1548 794 1552
rect 798 1548 802 1552
rect 910 1548 914 1552
rect 926 1548 930 1552
rect 942 1548 946 1552
rect 1022 1548 1026 1552
rect 1038 1548 1042 1552
rect 1062 1548 1066 1552
rect 1078 1548 1082 1552
rect 1094 1548 1098 1552
rect 1222 1558 1226 1562
rect 1254 1558 1258 1562
rect 1286 1558 1290 1562
rect 1158 1548 1162 1552
rect 1174 1548 1178 1552
rect 1230 1548 1234 1552
rect 1262 1548 1266 1552
rect 1366 1558 1370 1562
rect 1398 1558 1402 1562
rect 1446 1558 1450 1562
rect 1478 1558 1482 1562
rect 1526 1558 1530 1562
rect 1582 1558 1586 1562
rect 1766 1558 1770 1562
rect 1942 1558 1946 1562
rect 1998 1558 2002 1562
rect 2094 1558 2098 1562
rect 2190 1558 2194 1562
rect 1334 1548 1338 1552
rect 1342 1548 1346 1552
rect 1358 1548 1362 1552
rect 1398 1548 1402 1552
rect 1414 1548 1418 1552
rect 1462 1548 1466 1552
rect 1478 1548 1482 1552
rect 1558 1548 1562 1552
rect 1574 1548 1578 1552
rect 1598 1548 1602 1552
rect 1614 1548 1618 1552
rect 1694 1548 1698 1552
rect 1710 1548 1714 1552
rect 1726 1548 1730 1552
rect 1734 1548 1738 1552
rect 1798 1548 1802 1552
rect 1814 1548 1818 1552
rect 1846 1548 1850 1552
rect 1862 1548 1866 1552
rect 1894 1548 1898 1552
rect 1910 1548 1914 1552
rect 1958 1548 1962 1552
rect 1974 1548 1978 1552
rect 2014 1548 2018 1552
rect 2030 1548 2034 1552
rect 2078 1548 2082 1552
rect 2086 1548 2090 1552
rect 2118 1548 2122 1552
rect 2126 1548 2130 1552
rect 2134 1548 2138 1552
rect 2158 1548 2162 1552
rect 2262 1558 2266 1562
rect 2310 1558 2314 1562
rect 2382 1558 2386 1562
rect 2414 1558 2418 1562
rect 2510 1558 2514 1562
rect 2742 1558 2746 1562
rect 2838 1558 2842 1562
rect 2878 1558 2882 1562
rect 2894 1558 2898 1562
rect 2982 1558 2986 1562
rect 3142 1558 3146 1562
rect 3174 1558 3178 1562
rect 3334 1558 3338 1562
rect 3390 1558 3394 1562
rect 3422 1558 3426 1562
rect 3542 1558 3546 1562
rect 2214 1548 2218 1552
rect 2286 1548 2290 1552
rect 2374 1548 2378 1552
rect 2390 1548 2394 1552
rect 2398 1548 2402 1552
rect 2414 1548 2418 1552
rect 2502 1548 2506 1552
rect 2566 1548 2570 1552
rect 2598 1548 2602 1552
rect 2630 1548 2634 1552
rect 2654 1548 2658 1552
rect 2686 1548 2690 1552
rect 38 1538 42 1542
rect 54 1538 58 1542
rect 94 1538 98 1542
rect 118 1538 122 1542
rect 166 1538 170 1542
rect 174 1538 178 1542
rect 286 1538 290 1542
rect 294 1538 298 1542
rect 422 1538 426 1542
rect 454 1538 458 1542
rect 494 1538 498 1542
rect 542 1538 546 1542
rect 574 1538 578 1542
rect 606 1538 610 1542
rect 758 1538 762 1542
rect 806 1538 810 1542
rect 814 1538 818 1542
rect 830 1538 834 1542
rect 870 1538 874 1542
rect 934 1538 938 1542
rect 966 1538 970 1542
rect 1006 1538 1010 1542
rect 1030 1538 1034 1542
rect 1086 1538 1090 1542
rect 1110 1538 1114 1542
rect 1118 1538 1122 1542
rect 1166 1538 1170 1542
rect 1174 1538 1178 1542
rect 1206 1538 1210 1542
rect 1230 1538 1234 1542
rect 1262 1538 1266 1542
rect 1310 1538 1314 1542
rect 1318 1538 1322 1542
rect 1390 1538 1394 1542
rect 1414 1538 1418 1542
rect 1422 1538 1426 1542
rect 1454 1538 1458 1542
rect 1518 1538 1522 1542
rect 1542 1538 1546 1542
rect 1566 1538 1570 1542
rect 1606 1538 1610 1542
rect 1622 1538 1626 1542
rect 1630 1538 1634 1542
rect 1638 1538 1642 1542
rect 1654 1540 1658 1544
rect 1702 1538 1706 1542
rect 1718 1538 1722 1542
rect 1734 1538 1738 1542
rect 1750 1538 1754 1542
rect 1822 1538 1826 1542
rect 1838 1538 1842 1542
rect 1854 1538 1858 1542
rect 1870 1538 1874 1542
rect 1902 1538 1906 1542
rect 1918 1538 1922 1542
rect 1966 1538 1970 1542
rect 2022 1538 2026 1542
rect 2110 1538 2114 1542
rect 2174 1538 2178 1542
rect 2222 1538 2226 1542
rect 2230 1538 2234 1542
rect 2270 1538 2274 1542
rect 2286 1538 2290 1542
rect 2294 1538 2298 1542
rect 2318 1538 2322 1542
rect 2366 1538 2370 1542
rect 2406 1538 2410 1542
rect 2718 1548 2722 1552
rect 2750 1548 2754 1552
rect 2830 1548 2834 1552
rect 2854 1548 2858 1552
rect 2870 1548 2874 1552
rect 2950 1548 2954 1552
rect 2958 1548 2962 1552
rect 2990 1548 2994 1552
rect 3014 1548 3018 1552
rect 3030 1548 3034 1552
rect 3078 1548 3082 1552
rect 3118 1548 3122 1552
rect 3166 1548 3170 1552
rect 3206 1548 3210 1552
rect 3270 1548 3274 1552
rect 3286 1548 3290 1552
rect 3350 1548 3354 1552
rect 3366 1548 3370 1552
rect 3406 1548 3410 1552
rect 3438 1548 3442 1552
rect 3478 1548 3482 1552
rect 3486 1548 3490 1552
rect 3534 1548 3538 1552
rect 2430 1538 2434 1542
rect 2462 1538 2466 1542
rect 2526 1538 2530 1542
rect 2558 1538 2562 1542
rect 2606 1538 2610 1542
rect 2662 1538 2666 1542
rect 2678 1538 2682 1542
rect 2710 1538 2714 1542
rect 2790 1538 2794 1542
rect 2822 1538 2826 1542
rect 2862 1538 2866 1542
rect 2910 1538 2914 1542
rect 2926 1538 2930 1542
rect 2950 1538 2954 1542
rect 3126 1538 3130 1542
rect 3182 1538 3186 1542
rect 3214 1538 3218 1542
rect 3230 1538 3234 1542
rect 3366 1538 3370 1542
rect 3414 1538 3418 1542
rect 3446 1538 3450 1542
rect 3470 1538 3474 1542
rect 3526 1538 3530 1542
rect 3558 1538 3562 1542
rect 150 1528 154 1532
rect 262 1528 266 1532
rect 374 1528 378 1532
rect 566 1528 570 1532
rect 686 1528 690 1532
rect 694 1528 698 1532
rect 710 1528 714 1532
rect 838 1528 842 1532
rect 894 1528 898 1532
rect 958 1528 962 1532
rect 1278 1528 1282 1532
rect 1358 1528 1362 1532
rect 1486 1528 1490 1532
rect 1502 1528 1506 1532
rect 1550 1528 1554 1532
rect 1638 1528 1642 1532
rect 1678 1528 1682 1532
rect 1694 1528 1698 1532
rect 1766 1528 1770 1532
rect 1814 1528 1818 1532
rect 1886 1528 1890 1532
rect 1990 1528 1994 1532
rect 2094 1528 2098 1532
rect 2246 1528 2250 1532
rect 2318 1528 2322 1532
rect 2446 1528 2450 1532
rect 2454 1528 2458 1532
rect 2518 1528 2522 1532
rect 2582 1528 2586 1532
rect 2590 1528 2594 1532
rect 2622 1528 2626 1532
rect 2646 1528 2650 1532
rect 2678 1528 2682 1532
rect 2734 1528 2738 1532
rect 2798 1528 2802 1532
rect 2806 1528 2810 1532
rect 2886 1528 2890 1532
rect 2918 1528 2922 1532
rect 2926 1528 2930 1532
rect 2934 1528 2938 1532
rect 2974 1528 2978 1532
rect 3030 1528 3034 1532
rect 3070 1528 3074 1532
rect 3142 1528 3146 1532
rect 3230 1528 3234 1532
rect 3454 1528 3458 1532
rect 3510 1528 3514 1532
rect 46 1518 50 1522
rect 70 1518 74 1522
rect 182 1518 186 1522
rect 254 1518 258 1522
rect 270 1518 274 1522
rect 350 1518 354 1522
rect 382 1518 386 1522
rect 438 1518 442 1522
rect 470 1518 474 1522
rect 518 1518 522 1522
rect 598 1518 602 1522
rect 638 1518 642 1522
rect 702 1518 706 1522
rect 822 1518 826 1522
rect 862 1518 866 1522
rect 974 1518 978 1522
rect 1054 1518 1058 1522
rect 1062 1518 1066 1522
rect 1142 1518 1146 1522
rect 1198 1518 1202 1522
rect 1286 1518 1290 1522
rect 1334 1518 1338 1522
rect 1350 1518 1354 1522
rect 1518 1518 1522 1522
rect 1782 1518 1786 1522
rect 1982 1518 1986 1522
rect 2358 1518 2362 1522
rect 2614 1518 2618 1522
rect 2638 1518 2642 1522
rect 2670 1518 2674 1522
rect 2966 1518 2970 1522
rect 3022 1518 3026 1522
rect 3102 1518 3106 1522
rect 3222 1518 3226 1522
rect 3326 1518 3330 1522
rect 3462 1518 3466 1522
rect 994 1503 998 1507
rect 1001 1503 1005 1507
rect 2026 1503 2030 1507
rect 2033 1503 2037 1507
rect 3042 1503 3046 1507
rect 3049 1503 3053 1507
rect 446 1488 450 1492
rect 670 1488 674 1492
rect 702 1488 706 1492
rect 838 1488 842 1492
rect 1038 1488 1042 1492
rect 1134 1488 1138 1492
rect 1214 1488 1218 1492
rect 1366 1488 1370 1492
rect 1478 1488 1482 1492
rect 1534 1488 1538 1492
rect 1574 1488 1578 1492
rect 1590 1488 1594 1492
rect 1630 1488 1634 1492
rect 1686 1488 1690 1492
rect 1766 1488 1770 1492
rect 1862 1488 1866 1492
rect 1886 1488 1890 1492
rect 1934 1488 1938 1492
rect 1990 1488 1994 1492
rect 2046 1488 2050 1492
rect 2078 1488 2082 1492
rect 2102 1488 2106 1492
rect 2166 1488 2170 1492
rect 2318 1488 2322 1492
rect 2398 1488 2402 1492
rect 2534 1488 2538 1492
rect 2582 1488 2586 1492
rect 2622 1488 2626 1492
rect 2878 1488 2882 1492
rect 3166 1488 3170 1492
rect 3302 1488 3306 1492
rect 3382 1488 3386 1492
rect 3398 1488 3402 1492
rect 3518 1488 3522 1492
rect 6 1478 10 1482
rect 94 1478 98 1482
rect 326 1478 330 1482
rect 334 1478 338 1482
rect 350 1478 354 1482
rect 798 1478 802 1482
rect 846 1478 850 1482
rect 1270 1478 1274 1482
rect 1534 1478 1538 1482
rect 54 1468 58 1472
rect 102 1468 106 1472
rect 126 1468 130 1472
rect 174 1468 178 1472
rect 206 1468 210 1472
rect 286 1468 290 1472
rect 294 1468 298 1472
rect 382 1468 386 1472
rect 390 1468 394 1472
rect 422 1468 426 1472
rect 454 1468 458 1472
rect 486 1468 490 1472
rect 606 1468 610 1472
rect 654 1468 658 1472
rect 662 1468 666 1472
rect 710 1468 714 1472
rect 742 1468 746 1472
rect 774 1468 778 1472
rect 910 1468 914 1472
rect 918 1468 922 1472
rect 942 1468 946 1472
rect 974 1468 978 1472
rect 1182 1468 1186 1472
rect 1190 1468 1194 1472
rect 1222 1468 1226 1472
rect 1278 1468 1282 1472
rect 1302 1468 1306 1472
rect 1310 1468 1314 1472
rect 1342 1468 1346 1472
rect 1414 1468 1418 1472
rect 1470 1468 1474 1472
rect 1486 1468 1490 1472
rect 1494 1468 1498 1472
rect 1550 1468 1554 1472
rect 1558 1468 1562 1472
rect 1646 1478 1650 1482
rect 1662 1478 1666 1482
rect 1694 1478 1698 1482
rect 1726 1478 1730 1482
rect 1758 1478 1762 1482
rect 1790 1478 1794 1482
rect 1982 1478 1986 1482
rect 2094 1478 2098 1482
rect 2158 1478 2162 1482
rect 2286 1478 2290 1482
rect 2310 1478 2314 1482
rect 2366 1478 2370 1482
rect 2390 1478 2394 1482
rect 2558 1478 2562 1482
rect 2590 1478 2594 1482
rect 2686 1478 2690 1482
rect 2726 1478 2730 1482
rect 2758 1478 2762 1482
rect 2798 1478 2802 1482
rect 2822 1478 2826 1482
rect 2870 1478 2874 1482
rect 2902 1478 2906 1482
rect 2942 1478 2946 1482
rect 3014 1478 3018 1482
rect 3054 1478 3058 1482
rect 3270 1478 3274 1482
rect 3358 1478 3362 1482
rect 3390 1478 3394 1482
rect 3470 1478 3474 1482
rect 3510 1478 3514 1482
rect 1590 1468 1594 1472
rect 1606 1468 1610 1472
rect 1622 1468 1626 1472
rect 1678 1468 1682 1472
rect 1694 1468 1698 1472
rect 1742 1468 1746 1472
rect 1766 1468 1770 1472
rect 1782 1468 1786 1472
rect 1806 1468 1810 1472
rect 1838 1468 1842 1472
rect 1870 1468 1874 1472
rect 1878 1468 1882 1472
rect 1902 1468 1906 1472
rect 1958 1468 1962 1472
rect 2014 1468 2018 1472
rect 2086 1468 2090 1472
rect 2110 1468 2114 1472
rect 2126 1468 2130 1472
rect 2182 1468 2186 1472
rect 2206 1468 2210 1472
rect 2214 1468 2218 1472
rect 2406 1468 2410 1472
rect 2422 1468 2426 1472
rect 2438 1468 2442 1472
rect 2454 1468 2458 1472
rect 22 1458 26 1462
rect 102 1458 106 1462
rect 166 1458 170 1462
rect 198 1458 202 1462
rect 222 1458 226 1462
rect 246 1458 250 1462
rect 254 1458 258 1462
rect 278 1458 282 1462
rect 334 1458 338 1462
rect 374 1458 378 1462
rect 398 1458 402 1462
rect 446 1458 450 1462
rect 462 1458 466 1462
rect 478 1458 482 1462
rect 510 1458 514 1462
rect 542 1458 546 1462
rect 550 1458 554 1462
rect 566 1458 570 1462
rect 590 1458 594 1462
rect 598 1458 602 1462
rect 614 1458 618 1462
rect 686 1458 690 1462
rect 750 1458 754 1462
rect 766 1458 770 1462
rect 822 1458 826 1462
rect 870 1458 874 1462
rect 950 1458 954 1462
rect 974 1458 978 1462
rect 1014 1458 1018 1462
rect 1022 1458 1026 1462
rect 1062 1458 1066 1462
rect 1070 1458 1074 1462
rect 1094 1458 1098 1462
rect 1102 1458 1106 1462
rect 1110 1458 1114 1462
rect 1142 1458 1146 1462
rect 1150 1458 1154 1462
rect 1174 1458 1178 1462
rect 1198 1458 1202 1462
rect 1230 1458 1234 1462
rect 1254 1458 1258 1462
rect 1318 1458 1322 1462
rect 1342 1458 1346 1462
rect 1350 1458 1354 1462
rect 1374 1458 1378 1462
rect 1382 1458 1386 1462
rect 1406 1458 1410 1462
rect 1422 1458 1426 1462
rect 1430 1458 1434 1462
rect 1454 1458 1458 1462
rect 1486 1458 1490 1462
rect 1558 1458 1562 1462
rect 1614 1458 1618 1462
rect 1646 1458 1650 1462
rect 1670 1458 1674 1462
rect 1702 1458 1706 1462
rect 1734 1458 1738 1462
rect 1806 1458 1810 1462
rect 1862 1458 1866 1462
rect 1910 1458 1914 1462
rect 1950 1458 1954 1462
rect 1966 1458 1970 1462
rect 2006 1458 2010 1462
rect 2070 1458 2074 1462
rect 2118 1458 2122 1462
rect 2134 1458 2138 1462
rect 2150 1458 2154 1462
rect 2174 1458 2178 1462
rect 2198 1458 2202 1462
rect 2222 1458 2226 1462
rect 2238 1458 2242 1462
rect 2278 1458 2282 1462
rect 2310 1458 2314 1462
rect 2326 1458 2330 1462
rect 2358 1458 2362 1462
rect 2414 1458 2418 1462
rect 2430 1458 2434 1462
rect 2454 1458 2458 1462
rect 2486 1468 2490 1472
rect 2558 1468 2562 1472
rect 2598 1468 2602 1472
rect 2678 1468 2682 1472
rect 2742 1468 2746 1472
rect 2846 1468 2850 1472
rect 2862 1468 2866 1472
rect 2886 1468 2890 1472
rect 2958 1468 2962 1472
rect 2974 1468 2978 1472
rect 2982 1468 2986 1472
rect 3006 1468 3010 1472
rect 3022 1468 3026 1472
rect 3038 1468 3042 1472
rect 3070 1468 3074 1472
rect 3230 1468 3234 1472
rect 3238 1468 3242 1472
rect 3294 1468 3298 1472
rect 3326 1468 3330 1472
rect 3350 1468 3354 1472
rect 3366 1468 3370 1472
rect 3406 1468 3410 1472
rect 3430 1468 3434 1472
rect 3446 1468 3450 1472
rect 3454 1468 3458 1472
rect 3478 1468 3482 1472
rect 3526 1468 3530 1472
rect 3542 1468 3546 1472
rect 3558 1468 3562 1472
rect 2486 1458 2490 1462
rect 2518 1458 2522 1462
rect 2558 1458 2562 1462
rect 2606 1458 2610 1462
rect 2630 1458 2634 1462
rect 2662 1458 2666 1462
rect 2710 1458 2714 1462
rect 2766 1458 2770 1462
rect 2782 1458 2786 1462
rect 2838 1458 2842 1462
rect 2854 1458 2858 1462
rect 2902 1458 2906 1462
rect 2910 1458 2914 1462
rect 2918 1458 2922 1462
rect 2926 1458 2930 1462
rect 2950 1458 2954 1462
rect 2966 1458 2970 1462
rect 2990 1458 2994 1462
rect 3030 1458 3034 1462
rect 3102 1459 3106 1463
rect 3134 1458 3138 1462
rect 3174 1458 3178 1462
rect 3190 1458 3194 1462
rect 3230 1458 3234 1462
rect 3246 1458 3250 1462
rect 3270 1458 3274 1462
rect 3286 1458 3290 1462
rect 3318 1458 3322 1462
rect 3414 1458 3418 1462
rect 3438 1458 3442 1462
rect 3454 1458 3458 1462
rect 3502 1458 3506 1462
rect 46 1448 50 1452
rect 78 1448 82 1452
rect 94 1448 98 1452
rect 118 1448 122 1452
rect 142 1448 146 1452
rect 182 1448 186 1452
rect 262 1448 266 1452
rect 310 1448 314 1452
rect 358 1448 362 1452
rect 414 1448 418 1452
rect 462 1448 466 1452
rect 638 1448 642 1452
rect 678 1448 682 1452
rect 766 1448 770 1452
rect 790 1448 794 1452
rect 838 1448 842 1452
rect 894 1448 898 1452
rect 934 1448 938 1452
rect 1006 1448 1010 1452
rect 1158 1448 1162 1452
rect 1246 1448 1250 1452
rect 1286 1448 1290 1452
rect 1334 1448 1338 1452
rect 1366 1448 1370 1452
rect 1470 1448 1474 1452
rect 1518 1448 1522 1452
rect 1590 1448 1594 1452
rect 1766 1448 1770 1452
rect 1830 1448 1834 1452
rect 1894 1448 1898 1452
rect 1926 1448 1930 1452
rect 1934 1448 1938 1452
rect 1990 1448 1994 1452
rect 2070 1448 2074 1452
rect 2150 1448 2154 1452
rect 2182 1448 2186 1452
rect 2238 1448 2242 1452
rect 2462 1448 2466 1452
rect 2470 1448 2474 1452
rect 2510 1448 2514 1452
rect 2662 1448 2666 1452
rect 2678 1448 2682 1452
rect 2726 1448 2730 1452
rect 2766 1448 2770 1452
rect 2838 1448 2842 1452
rect 2990 1448 2994 1452
rect 3174 1448 3178 1452
rect 3206 1448 3210 1452
rect 3222 1448 3226 1452
rect 3270 1448 3274 1452
rect 3326 1448 3330 1452
rect 3382 1448 3386 1452
rect 3422 1448 3426 1452
rect 3542 1448 3546 1452
rect 238 1438 242 1442
rect 614 1438 618 1442
rect 870 1438 874 1442
rect 918 1438 922 1442
rect 1726 1438 1730 1442
rect 1790 1438 1794 1442
rect 2254 1438 2258 1442
rect 3022 1438 3026 1442
rect 62 1428 66 1432
rect 782 1428 786 1432
rect 1086 1428 1090 1432
rect 1174 1428 1178 1432
rect 30 1418 34 1422
rect 86 1418 90 1422
rect 166 1418 170 1422
rect 198 1418 202 1422
rect 278 1418 282 1422
rect 302 1418 306 1422
rect 318 1418 322 1422
rect 374 1418 378 1422
rect 534 1418 538 1422
rect 582 1418 586 1422
rect 726 1418 730 1422
rect 1398 1418 1402 1422
rect 1646 1418 1650 1422
rect 1910 1418 1914 1422
rect 1950 1418 1954 1422
rect 1974 1418 1978 1422
rect 2342 1418 2346 1422
rect 2374 1418 2378 1422
rect 2782 1418 2786 1422
rect 2926 1418 2930 1422
rect 3054 1418 3058 1422
rect 482 1403 486 1407
rect 489 1403 493 1407
rect 1514 1403 1518 1407
rect 1521 1403 1525 1407
rect 2538 1403 2542 1407
rect 2545 1403 2549 1407
rect 510 1388 514 1392
rect 814 1388 818 1392
rect 894 1388 898 1392
rect 942 1388 946 1392
rect 1278 1388 1282 1392
rect 1310 1388 1314 1392
rect 1382 1388 1386 1392
rect 1446 1388 1450 1392
rect 1678 1388 1682 1392
rect 1742 1388 1746 1392
rect 1782 1388 1786 1392
rect 1918 1388 1922 1392
rect 2254 1388 2258 1392
rect 2270 1388 2274 1392
rect 2414 1388 2418 1392
rect 2510 1388 2514 1392
rect 2862 1388 2866 1392
rect 2910 1388 2914 1392
rect 3062 1388 3066 1392
rect 3102 1388 3106 1392
rect 3150 1388 3154 1392
rect 3318 1388 3322 1392
rect 3398 1388 3402 1392
rect 3454 1388 3458 1392
rect 3542 1388 3546 1392
rect 2894 1378 2898 1382
rect 2990 1378 2994 1382
rect 606 1368 610 1372
rect 1734 1368 1738 1372
rect 2118 1368 2122 1372
rect 2510 1368 2514 1372
rect 2622 1368 2626 1372
rect 3278 1368 3282 1372
rect 3494 1368 3498 1372
rect 6 1358 10 1362
rect 30 1358 34 1362
rect 54 1358 58 1362
rect 102 1358 106 1362
rect 166 1358 170 1362
rect 182 1358 186 1362
rect 214 1358 218 1362
rect 230 1358 234 1362
rect 238 1358 242 1362
rect 310 1358 314 1362
rect 342 1358 346 1362
rect 350 1358 354 1362
rect 390 1358 394 1362
rect 398 1358 402 1362
rect 422 1358 426 1362
rect 470 1358 474 1362
rect 486 1358 490 1362
rect 574 1358 578 1362
rect 646 1358 650 1362
rect 670 1358 674 1362
rect 702 1358 706 1362
rect 734 1358 738 1362
rect 758 1358 762 1362
rect 782 1358 786 1362
rect 878 1358 882 1362
rect 902 1358 906 1362
rect 974 1358 978 1362
rect 982 1358 986 1362
rect 1030 1358 1034 1362
rect 1222 1358 1226 1362
rect 1238 1358 1242 1362
rect 1294 1358 1298 1362
rect 1326 1358 1330 1362
rect 1430 1358 1434 1362
rect 1462 1358 1466 1362
rect 1478 1358 1482 1362
rect 1494 1358 1498 1362
rect 1502 1358 1506 1362
rect 1526 1358 1530 1362
rect 1542 1358 1546 1362
rect 1558 1358 1562 1362
rect 1646 1358 1650 1362
rect 1734 1358 1738 1362
rect 1822 1358 1826 1362
rect 1830 1358 1834 1362
rect 1878 1358 1882 1362
rect 1902 1358 1906 1362
rect 1974 1358 1978 1362
rect 2102 1358 2106 1362
rect 2190 1358 2194 1362
rect 2222 1358 2226 1362
rect 2342 1358 2346 1362
rect 2502 1358 2506 1362
rect 2550 1358 2554 1362
rect 2606 1358 2610 1362
rect 2678 1358 2682 1362
rect 2686 1358 2690 1362
rect 2726 1358 2730 1362
rect 2782 1358 2786 1362
rect 2846 1358 2850 1362
rect 2966 1358 2970 1362
rect 2974 1358 2978 1362
rect 70 1348 74 1352
rect 86 1348 90 1352
rect 110 1348 114 1352
rect 254 1348 258 1352
rect 294 1348 298 1352
rect 326 1348 330 1352
rect 438 1348 442 1352
rect 454 1348 458 1352
rect 526 1348 530 1352
rect 534 1348 538 1352
rect 558 1348 562 1352
rect 606 1348 610 1352
rect 686 1348 690 1352
rect 718 1348 722 1352
rect 734 1348 738 1352
rect 790 1348 794 1352
rect 798 1348 802 1352
rect 830 1348 834 1352
rect 862 1348 866 1352
rect 926 1348 930 1352
rect 998 1348 1002 1352
rect 1054 1348 1058 1352
rect 1062 1348 1066 1352
rect 1086 1348 1090 1352
rect 1102 1348 1106 1352
rect 1134 1348 1138 1352
rect 1182 1348 1186 1352
rect 1214 1348 1218 1352
rect 1222 1348 1226 1352
rect 1246 1348 1250 1352
rect 1294 1348 1298 1352
rect 1310 1348 1314 1352
rect 1334 1348 1338 1352
rect 1350 1348 1354 1352
rect 1358 1348 1362 1352
rect 1366 1348 1370 1352
rect 1390 1348 1394 1352
rect 1414 1348 1418 1352
rect 1478 1348 1482 1352
rect 1566 1348 1570 1352
rect 1582 1348 1586 1352
rect 1590 1348 1594 1352
rect 1654 1348 1658 1352
rect 1662 1348 1666 1352
rect 1686 1348 1690 1352
rect 1726 1348 1730 1352
rect 1742 1348 1746 1352
rect 1766 1348 1770 1352
rect 1798 1348 1802 1352
rect 1814 1348 1818 1352
rect 1846 1348 1850 1352
rect 1910 1348 1914 1352
rect 1942 1348 1946 1352
rect 1958 1348 1962 1352
rect 1982 1348 1986 1352
rect 2054 1348 2058 1352
rect 22 1338 26 1342
rect 46 1338 50 1342
rect 86 1338 90 1342
rect 134 1338 138 1342
rect 142 1338 146 1342
rect 166 1338 170 1342
rect 190 1338 194 1342
rect 214 1338 218 1342
rect 246 1338 250 1342
rect 262 1338 266 1342
rect 318 1338 322 1342
rect 374 1338 378 1342
rect 414 1338 418 1342
rect 438 1338 442 1342
rect 446 1338 450 1342
rect 518 1338 522 1342
rect 590 1338 594 1342
rect 630 1338 634 1342
rect 646 1338 650 1342
rect 670 1338 674 1342
rect 710 1338 714 1342
rect 742 1338 746 1342
rect 758 1338 762 1342
rect 918 1338 922 1342
rect 958 1338 962 1342
rect 990 1338 994 1342
rect 1006 1338 1010 1342
rect 1046 1338 1050 1342
rect 1102 1338 1106 1342
rect 1110 1338 1114 1342
rect 1174 1338 1178 1342
rect 1214 1338 1218 1342
rect 1270 1338 1274 1342
rect 2094 1348 2098 1352
rect 2110 1348 2114 1352
rect 2158 1348 2162 1352
rect 2174 1348 2178 1352
rect 2206 1348 2210 1352
rect 2230 1348 2234 1352
rect 2270 1348 2274 1352
rect 2294 1348 2298 1352
rect 2318 1348 2322 1352
rect 2358 1348 2362 1352
rect 2430 1348 2434 1352
rect 1406 1338 1410 1342
rect 1438 1338 1442 1342
rect 1470 1338 1474 1342
rect 1518 1338 1522 1342
rect 1542 1338 1546 1342
rect 1558 1338 1562 1342
rect 1590 1338 1594 1342
rect 1622 1338 1626 1342
rect 1702 1338 1706 1342
rect 1790 1338 1794 1342
rect 1854 1338 1858 1342
rect 1902 1338 1906 1342
rect 1918 1338 1922 1342
rect 1934 1338 1938 1342
rect 1942 1338 1946 1342
rect 1990 1338 1994 1342
rect 2046 1338 2050 1342
rect 2062 1338 2066 1342
rect 2070 1338 2074 1342
rect 2086 1338 2090 1342
rect 2150 1338 2154 1342
rect 2166 1338 2170 1342
rect 2198 1338 2202 1342
rect 2214 1338 2218 1342
rect 2230 1338 2234 1342
rect 2262 1338 2266 1342
rect 2366 1338 2370 1342
rect 2390 1338 2394 1342
rect 2406 1338 2410 1342
rect 2478 1348 2482 1352
rect 2518 1348 2522 1352
rect 2566 1348 2570 1352
rect 2582 1348 2586 1352
rect 2614 1348 2618 1352
rect 2646 1348 2650 1352
rect 2654 1348 2658 1352
rect 2694 1348 2698 1352
rect 2702 1348 2706 1352
rect 2718 1348 2722 1352
rect 2750 1348 2754 1352
rect 2766 1348 2770 1352
rect 2814 1348 2818 1352
rect 2830 1348 2834 1352
rect 2870 1348 2874 1352
rect 2878 1348 2882 1352
rect 2926 1348 2930 1352
rect 2950 1348 2954 1352
rect 2990 1348 2994 1352
rect 3006 1348 3010 1352
rect 3030 1348 3034 1352
rect 3078 1348 3082 1352
rect 3086 1348 3090 1352
rect 3206 1358 3210 1362
rect 3350 1358 3354 1362
rect 3438 1358 3442 1362
rect 3526 1358 3530 1362
rect 3534 1358 3538 1362
rect 3222 1348 3226 1352
rect 3238 1348 3242 1352
rect 3278 1348 3282 1352
rect 3286 1348 3290 1352
rect 3342 1348 3346 1352
rect 3366 1348 3370 1352
rect 3454 1348 3458 1352
rect 3470 1348 3474 1352
rect 3510 1348 3514 1352
rect 3534 1348 3538 1352
rect 2574 1338 2578 1342
rect 2582 1338 2586 1342
rect 2622 1338 2626 1342
rect 2638 1338 2642 1342
rect 2654 1338 2658 1342
rect 2710 1338 2714 1342
rect 2726 1338 2730 1342
rect 2742 1338 2746 1342
rect 2758 1338 2762 1342
rect 2806 1338 2810 1342
rect 2822 1338 2826 1342
rect 2934 1338 2938 1342
rect 2942 1338 2946 1342
rect 2958 1338 2962 1342
rect 2998 1338 3002 1342
rect 3118 1338 3122 1342
rect 3166 1338 3170 1342
rect 3174 1338 3178 1342
rect 3190 1338 3194 1342
rect 3230 1338 3234 1342
rect 3334 1338 3338 1342
rect 3358 1338 3362 1342
rect 3374 1338 3378 1342
rect 3382 1338 3386 1342
rect 3462 1338 3466 1342
rect 3478 1338 3482 1342
rect 3502 1338 3506 1342
rect 3550 1338 3554 1342
rect 270 1328 274 1332
rect 310 1328 314 1332
rect 838 1328 842 1332
rect 886 1328 890 1332
rect 1126 1328 1130 1332
rect 1150 1328 1154 1332
rect 1190 1328 1194 1332
rect 1262 1328 1266 1332
rect 1350 1328 1354 1332
rect 1566 1328 1570 1332
rect 1614 1328 1618 1332
rect 1838 1328 1842 1332
rect 1878 1328 1882 1332
rect 2014 1328 2018 1332
rect 2134 1328 2138 1332
rect 2190 1328 2194 1332
rect 2254 1328 2258 1332
rect 2334 1328 2338 1332
rect 2374 1328 2378 1332
rect 2446 1328 2450 1332
rect 2470 1328 2474 1332
rect 2494 1328 2498 1332
rect 2678 1328 2682 1332
rect 2846 1328 2850 1332
rect 2854 1328 2858 1332
rect 3254 1328 3258 1332
rect 3318 1328 3322 1332
rect 3494 1328 3498 1332
rect 14 1318 18 1322
rect 38 1318 42 1322
rect 54 1318 58 1322
rect 94 1318 98 1322
rect 150 1318 154 1322
rect 174 1318 178 1322
rect 206 1318 210 1322
rect 230 1318 234 1322
rect 342 1318 346 1322
rect 350 1318 354 1322
rect 382 1318 386 1322
rect 398 1318 402 1322
rect 486 1318 490 1322
rect 550 1318 554 1322
rect 582 1318 586 1322
rect 670 1318 674 1322
rect 702 1318 706 1322
rect 734 1318 738 1322
rect 774 1318 778 1322
rect 878 1318 882 1322
rect 902 1318 906 1322
rect 966 1318 970 1322
rect 1038 1318 1042 1322
rect 1118 1318 1122 1322
rect 1166 1318 1170 1322
rect 1198 1318 1202 1322
rect 1646 1318 1650 1322
rect 1998 1318 2002 1322
rect 2038 1318 2042 1322
rect 2078 1318 2082 1322
rect 2110 1318 2114 1322
rect 2142 1318 2146 1322
rect 2342 1318 2346 1322
rect 2382 1318 2386 1322
rect 2534 1318 2538 1322
rect 2606 1318 2610 1322
rect 2798 1318 2802 1322
rect 3302 1318 3306 1322
rect 994 1303 998 1307
rect 1001 1303 1005 1307
rect 2026 1303 2030 1307
rect 2033 1303 2037 1307
rect 3042 1303 3046 1307
rect 3049 1303 3053 1307
rect 14 1288 18 1292
rect 62 1288 66 1292
rect 254 1288 258 1292
rect 366 1288 370 1292
rect 638 1288 642 1292
rect 702 1288 706 1292
rect 854 1288 858 1292
rect 886 1288 890 1292
rect 1094 1288 1098 1292
rect 1110 1288 1114 1292
rect 1222 1288 1226 1292
rect 1270 1288 1274 1292
rect 1294 1288 1298 1292
rect 1326 1288 1330 1292
rect 1382 1288 1386 1292
rect 1406 1288 1410 1292
rect 1438 1288 1442 1292
rect 1694 1288 1698 1292
rect 1854 1288 1858 1292
rect 1894 1288 1898 1292
rect 2102 1288 2106 1292
rect 2198 1288 2202 1292
rect 2238 1288 2242 1292
rect 2262 1288 2266 1292
rect 2302 1288 2306 1292
rect 2374 1288 2378 1292
rect 2430 1288 2434 1292
rect 2510 1288 2514 1292
rect 2558 1288 2562 1292
rect 2790 1288 2794 1292
rect 2846 1288 2850 1292
rect 2942 1288 2946 1292
rect 2990 1288 2994 1292
rect 3014 1288 3018 1292
rect 3086 1288 3090 1292
rect 3214 1288 3218 1292
rect 3430 1288 3434 1292
rect 3558 1288 3562 1292
rect 126 1278 130 1282
rect 166 1278 170 1282
rect 246 1278 250 1282
rect 446 1278 450 1282
rect 630 1278 634 1282
rect 710 1278 714 1282
rect 742 1278 746 1282
rect 846 1278 850 1282
rect 894 1278 898 1282
rect 998 1278 1002 1282
rect 1014 1278 1018 1282
rect 1022 1278 1026 1282
rect 1038 1278 1042 1282
rect 1046 1278 1050 1282
rect 158 1268 162 1272
rect 182 1268 186 1272
rect 198 1268 202 1272
rect 286 1268 290 1272
rect 302 1268 306 1272
rect 342 1268 346 1272
rect 430 1268 434 1272
rect 438 1268 442 1272
rect 526 1268 530 1272
rect 558 1268 562 1272
rect 590 1268 594 1272
rect 614 1268 618 1272
rect 662 1268 666 1272
rect 694 1268 698 1272
rect 726 1268 730 1272
rect 790 1268 794 1272
rect 806 1268 810 1272
rect 822 1268 826 1272
rect 830 1268 834 1272
rect 870 1268 874 1272
rect 926 1268 930 1272
rect 1022 1268 1026 1272
rect 1070 1268 1074 1272
rect 30 1258 34 1262
rect 46 1258 50 1262
rect 70 1258 74 1262
rect 78 1258 82 1262
rect 110 1258 114 1262
rect 134 1258 138 1262
rect 182 1258 186 1262
rect 214 1258 218 1262
rect 222 1258 226 1262
rect 270 1258 274 1262
rect 318 1258 322 1262
rect 350 1258 354 1262
rect 374 1258 378 1262
rect 398 1258 402 1262
rect 422 1258 426 1262
rect 454 1258 458 1262
rect 494 1258 498 1262
rect 502 1258 506 1262
rect 550 1258 554 1262
rect 566 1258 570 1262
rect 606 1258 610 1262
rect 654 1258 658 1262
rect 686 1258 690 1262
rect 718 1258 722 1262
rect 782 1258 786 1262
rect 814 1258 818 1262
rect 878 1258 882 1262
rect 942 1258 946 1262
rect 966 1258 970 1262
rect 974 1258 978 1262
rect 982 1258 986 1262
rect 1006 1258 1010 1262
rect 1062 1258 1066 1262
rect 1078 1258 1082 1262
rect 1102 1258 1106 1262
rect 1150 1278 1154 1282
rect 1206 1278 1210 1282
rect 1214 1278 1218 1282
rect 1262 1278 1266 1282
rect 1414 1278 1418 1282
rect 1462 1278 1466 1282
rect 1494 1278 1498 1282
rect 1574 1278 1578 1282
rect 1590 1278 1594 1282
rect 1686 1278 1690 1282
rect 1742 1278 1746 1282
rect 1750 1278 1754 1282
rect 1766 1278 1770 1282
rect 1966 1278 1970 1282
rect 1974 1278 1978 1282
rect 2038 1278 2042 1282
rect 2086 1278 2090 1282
rect 2094 1278 2098 1282
rect 2294 1278 2298 1282
rect 2350 1278 2354 1282
rect 2406 1278 2410 1282
rect 2438 1278 2442 1282
rect 2462 1278 2466 1282
rect 2486 1278 2490 1282
rect 2518 1278 2522 1282
rect 2582 1278 2586 1282
rect 2830 1278 2834 1282
rect 2894 1278 2898 1282
rect 2998 1278 3002 1282
rect 3150 1278 3154 1282
rect 3198 1278 3202 1282
rect 3254 1278 3258 1282
rect 1134 1268 1138 1272
rect 1150 1268 1154 1272
rect 1174 1268 1178 1272
rect 1254 1268 1258 1272
rect 1286 1268 1290 1272
rect 1318 1268 1322 1272
rect 1350 1268 1354 1272
rect 1390 1268 1394 1272
rect 1430 1268 1434 1272
rect 1446 1268 1450 1272
rect 1510 1268 1514 1272
rect 1542 1268 1546 1272
rect 1566 1268 1570 1272
rect 1598 1268 1602 1272
rect 1646 1268 1650 1272
rect 1126 1258 1130 1262
rect 1142 1258 1146 1262
rect 1182 1258 1186 1262
rect 1246 1258 1250 1262
rect 1278 1258 1282 1262
rect 1294 1258 1298 1262
rect 1310 1258 1314 1262
rect 1342 1258 1346 1262
rect 1350 1260 1354 1264
rect 1366 1258 1370 1262
rect 1390 1258 1394 1262
rect 1422 1258 1426 1262
rect 1454 1258 1458 1262
rect 1542 1258 1546 1262
rect 1574 1258 1578 1262
rect 1638 1258 1642 1262
rect 1646 1258 1650 1262
rect 1670 1268 1674 1272
rect 1702 1268 1706 1272
rect 1726 1268 1730 1272
rect 1790 1268 1794 1272
rect 1822 1268 1826 1272
rect 1830 1268 1834 1272
rect 1846 1268 1850 1272
rect 1878 1268 1882 1272
rect 1910 1268 1914 1272
rect 2006 1268 2010 1272
rect 2022 1268 2026 1272
rect 2110 1268 2114 1272
rect 2126 1268 2130 1272
rect 2206 1268 2210 1272
rect 2214 1268 2218 1272
rect 2246 1268 2250 1272
rect 2294 1268 2298 1272
rect 2310 1268 2314 1272
rect 2334 1268 2338 1272
rect 2390 1268 2394 1272
rect 2422 1268 2426 1272
rect 2502 1268 2506 1272
rect 2526 1268 2530 1272
rect 2542 1268 2546 1272
rect 2614 1268 2618 1272
rect 2654 1268 2658 1272
rect 2670 1268 2674 1272
rect 2694 1268 2698 1272
rect 2758 1268 2762 1272
rect 2854 1268 2858 1272
rect 2886 1268 2890 1272
rect 2918 1268 2922 1272
rect 2966 1268 2970 1272
rect 2974 1268 2978 1272
rect 3014 1268 3018 1272
rect 3030 1268 3034 1272
rect 3054 1268 3058 1272
rect 3102 1268 3106 1272
rect 3158 1268 3162 1272
rect 3206 1268 3210 1272
rect 3238 1268 3242 1272
rect 3278 1268 3282 1272
rect 3294 1268 3298 1272
rect 3422 1278 3426 1282
rect 3462 1278 3466 1282
rect 3310 1268 3314 1272
rect 3366 1268 3370 1272
rect 3398 1268 3402 1272
rect 3414 1268 3418 1272
rect 3478 1268 3482 1272
rect 1662 1258 1666 1262
rect 1710 1258 1714 1262
rect 1718 1258 1722 1262
rect 1766 1258 1770 1262
rect 1814 1258 1818 1262
rect 1870 1258 1874 1262
rect 1902 1258 1906 1262
rect 1918 1258 1922 1262
rect 1934 1258 1938 1262
rect 1950 1258 1954 1262
rect 1998 1258 2002 1262
rect 2070 1258 2074 1262
rect 2118 1258 2122 1262
rect 2134 1258 2138 1262
rect 2158 1258 2162 1262
rect 2190 1258 2194 1262
rect 2206 1258 2210 1262
rect 2318 1258 2322 1262
rect 2326 1258 2330 1262
rect 2382 1258 2386 1262
rect 2414 1258 2418 1262
rect 2446 1258 2450 1262
rect 2470 1258 2474 1262
rect 2494 1258 2498 1262
rect 2550 1258 2554 1262
rect 2582 1258 2586 1262
rect 2606 1258 2610 1262
rect 2630 1258 2634 1262
rect 2718 1258 2722 1262
rect 2734 1258 2738 1262
rect 2782 1258 2786 1262
rect 2814 1258 2818 1262
rect 2886 1258 2890 1262
rect 2894 1258 2898 1262
rect 2910 1258 2914 1262
rect 2926 1258 2930 1262
rect 3110 1258 3114 1262
rect 3166 1258 3170 1262
rect 3190 1258 3194 1262
rect 3238 1258 3242 1262
rect 3270 1258 3274 1262
rect 3350 1258 3354 1262
rect 3374 1258 3378 1262
rect 3438 1258 3442 1262
rect 3446 1258 3450 1262
rect 3494 1259 3498 1263
rect 86 1248 90 1252
rect 182 1248 186 1252
rect 198 1248 202 1252
rect 230 1248 234 1252
rect 254 1248 258 1252
rect 294 1248 298 1252
rect 302 1248 306 1252
rect 334 1248 338 1252
rect 366 1248 370 1252
rect 406 1248 410 1252
rect 454 1248 458 1252
rect 478 1248 482 1252
rect 582 1248 586 1252
rect 590 1248 594 1252
rect 638 1248 642 1252
rect 670 1248 674 1252
rect 798 1248 802 1252
rect 854 1248 858 1252
rect 902 1248 906 1252
rect 918 1248 922 1252
rect 1094 1248 1098 1252
rect 1174 1248 1178 1252
rect 1230 1248 1234 1252
rect 1326 1248 1330 1252
rect 1502 1248 1506 1252
rect 1534 1248 1538 1252
rect 1550 1248 1554 1252
rect 1614 1248 1618 1252
rect 1678 1248 1682 1252
rect 1774 1248 1778 1252
rect 1846 1248 1850 1252
rect 1886 1248 1890 1252
rect 1934 1248 1938 1252
rect 2006 1248 2010 1252
rect 2150 1248 2154 1252
rect 2158 1248 2162 1252
rect 2190 1248 2194 1252
rect 2238 1248 2242 1252
rect 2262 1248 2266 1252
rect 2286 1248 2290 1252
rect 2374 1248 2378 1252
rect 2478 1248 2482 1252
rect 2542 1248 2546 1252
rect 2590 1248 2594 1252
rect 2622 1248 2626 1252
rect 2726 1248 2730 1252
rect 2774 1248 2778 1252
rect 2838 1248 2842 1252
rect 2862 1248 2866 1252
rect 2878 1248 2882 1252
rect 2942 1248 2946 1252
rect 2950 1248 2954 1252
rect 3014 1248 3018 1252
rect 3126 1248 3130 1252
rect 3182 1248 3186 1252
rect 3206 1248 3210 1252
rect 3278 1248 3282 1252
rect 3294 1248 3298 1252
rect 3358 1248 3362 1252
rect 3398 1248 3402 1252
rect 246 1238 250 1242
rect 422 1238 426 1242
rect 598 1238 602 1242
rect 1062 1238 1066 1242
rect 1246 1238 1250 1242
rect 1566 1238 1570 1242
rect 2638 1238 2642 1242
rect 2742 1238 2746 1242
rect 3342 1238 3346 1242
rect 1166 1228 1170 1232
rect 1742 1228 1746 1232
rect 1814 1228 1818 1232
rect 2038 1228 2042 1232
rect 3326 1228 3330 1232
rect 102 1218 106 1222
rect 318 1218 322 1222
rect 534 1218 538 1222
rect 686 1218 690 1222
rect 742 1218 746 1222
rect 782 1218 786 1222
rect 958 1218 962 1222
rect 1206 1218 1210 1222
rect 1638 1218 1642 1222
rect 1974 1218 1978 1222
rect 2014 1218 2018 1222
rect 2174 1218 2178 1222
rect 2406 1218 2410 1222
rect 2446 1218 2450 1222
rect 2646 1218 2650 1222
rect 2662 1218 2666 1222
rect 2750 1218 2754 1222
rect 3350 1218 3354 1222
rect 3446 1218 3450 1222
rect 482 1203 486 1207
rect 489 1203 493 1207
rect 1514 1203 1518 1207
rect 1521 1203 1525 1207
rect 2538 1203 2542 1207
rect 2545 1203 2549 1207
rect 14 1188 18 1192
rect 142 1188 146 1192
rect 238 1188 242 1192
rect 342 1188 346 1192
rect 502 1188 506 1192
rect 566 1188 570 1192
rect 1022 1188 1026 1192
rect 1078 1188 1082 1192
rect 1278 1188 1282 1192
rect 1310 1188 1314 1192
rect 1438 1188 1442 1192
rect 1558 1188 1562 1192
rect 1638 1188 1642 1192
rect 1734 1188 1738 1192
rect 1790 1188 1794 1192
rect 1862 1188 1866 1192
rect 2022 1188 2026 1192
rect 2062 1188 2066 1192
rect 2126 1188 2130 1192
rect 2214 1188 2218 1192
rect 2342 1188 2346 1192
rect 2558 1188 2562 1192
rect 2574 1188 2578 1192
rect 2918 1188 2922 1192
rect 2942 1188 2946 1192
rect 2966 1188 2970 1192
rect 3014 1188 3018 1192
rect 3070 1188 3074 1192
rect 3406 1188 3410 1192
rect 398 1178 402 1182
rect 1350 1178 1354 1182
rect 2870 1178 2874 1182
rect 3558 1178 3562 1182
rect 294 1168 298 1172
rect 1158 1168 1162 1172
rect 1470 1168 1474 1172
rect 1902 1168 1906 1172
rect 3398 1168 3402 1172
rect 3406 1168 3410 1172
rect 3526 1168 3530 1172
rect 30 1158 34 1162
rect 62 1158 66 1162
rect 86 1158 90 1162
rect 126 1158 130 1162
rect 158 1158 162 1162
rect 166 1158 170 1162
rect 182 1158 186 1162
rect 222 1158 226 1162
rect 318 1158 322 1162
rect 358 1158 362 1162
rect 414 1158 418 1162
rect 446 1158 450 1162
rect 550 1158 554 1162
rect 582 1158 586 1162
rect 654 1158 658 1162
rect 14 1148 18 1152
rect 30 1148 34 1152
rect 142 1148 146 1152
rect 190 1148 194 1152
rect 206 1148 210 1152
rect 238 1148 242 1152
rect 278 1148 282 1152
rect 302 1148 306 1152
rect 310 1148 314 1152
rect 374 1148 378 1152
rect 398 1148 402 1152
rect 446 1148 450 1152
rect 470 1148 474 1152
rect 518 1148 522 1152
rect 534 1148 538 1152
rect 558 1148 562 1152
rect 614 1148 618 1152
rect 638 1148 642 1152
rect 646 1148 650 1152
rect 686 1148 690 1152
rect 718 1148 722 1152
rect 742 1148 746 1152
rect 750 1148 754 1152
rect 766 1148 770 1152
rect 790 1158 794 1162
rect 814 1158 818 1162
rect 870 1158 874 1162
rect 966 1158 970 1162
rect 990 1158 994 1162
rect 1038 1158 1042 1162
rect 1062 1158 1066 1162
rect 1190 1158 1194 1162
rect 1206 1158 1210 1162
rect 1254 1158 1258 1162
rect 830 1148 834 1152
rect 846 1148 850 1152
rect 878 1148 882 1152
rect 6 1138 10 1142
rect 38 1138 42 1142
rect 54 1138 58 1142
rect 70 1138 74 1142
rect 102 1138 106 1142
rect 110 1138 114 1142
rect 134 1138 138 1142
rect 182 1138 186 1142
rect 214 1138 218 1142
rect 334 1138 338 1142
rect 390 1138 394 1142
rect 422 1138 426 1142
rect 462 1138 466 1142
rect 534 1138 538 1142
rect 606 1138 610 1142
rect 662 1138 666 1142
rect 678 1138 682 1142
rect 686 1138 690 1142
rect 702 1138 706 1142
rect 758 1138 762 1142
rect 806 1138 810 1142
rect 822 1138 826 1142
rect 838 1138 842 1142
rect 846 1138 850 1142
rect 910 1148 914 1152
rect 934 1148 938 1152
rect 942 1148 946 1152
rect 1022 1148 1026 1152
rect 1038 1148 1042 1152
rect 1078 1148 1082 1152
rect 1086 1148 1090 1152
rect 1126 1148 1130 1152
rect 1134 1148 1138 1152
rect 1150 1148 1154 1152
rect 1174 1148 1178 1152
rect 1182 1148 1186 1152
rect 1206 1148 1210 1152
rect 1238 1148 1242 1152
rect 1390 1158 1394 1162
rect 1422 1158 1426 1162
rect 1454 1158 1458 1162
rect 1574 1158 1578 1162
rect 1654 1158 1658 1162
rect 1694 1158 1698 1162
rect 1766 1158 1770 1162
rect 1822 1158 1826 1162
rect 1830 1158 1834 1162
rect 2006 1158 2010 1162
rect 2038 1158 2042 1162
rect 2310 1158 2314 1162
rect 2742 1158 2746 1162
rect 2846 1158 2850 1162
rect 1278 1148 1282 1152
rect 1294 1148 1298 1152
rect 1302 1148 1306 1152
rect 1342 1148 1346 1152
rect 1350 1148 1354 1152
rect 1398 1148 1402 1152
rect 1438 1148 1442 1152
rect 1470 1148 1474 1152
rect 1486 1148 1490 1152
rect 1494 1148 1498 1152
rect 1518 1148 1522 1152
rect 1550 1148 1554 1152
rect 1558 1148 1562 1152
rect 1582 1148 1586 1152
rect 1590 1148 1594 1152
rect 1614 1148 1618 1152
rect 1638 1148 1642 1152
rect 1654 1148 1658 1152
rect 1678 1148 1682 1152
rect 1686 1148 1690 1152
rect 1734 1148 1738 1152
rect 1750 1148 1754 1152
rect 1774 1148 1778 1152
rect 1854 1148 1858 1152
rect 1870 1148 1874 1152
rect 1910 1148 1914 1152
rect 1934 1148 1938 1152
rect 1950 1148 1954 1152
rect 1966 1148 1970 1152
rect 1990 1148 1994 1152
rect 2078 1148 2082 1152
rect 2134 1148 2138 1152
rect 2174 1148 2178 1152
rect 2190 1148 2194 1152
rect 2206 1148 2210 1152
rect 2278 1148 2282 1152
rect 2374 1148 2378 1152
rect 2382 1148 2386 1152
rect 2414 1148 2418 1152
rect 2510 1148 2514 1152
rect 2518 1148 2522 1152
rect 2582 1148 2586 1152
rect 2614 1148 2618 1152
rect 2646 1148 2650 1152
rect 2678 1148 2682 1152
rect 2710 1148 2714 1152
rect 2726 1148 2730 1152
rect 2766 1148 2770 1152
rect 2782 1148 2786 1152
rect 2798 1148 2802 1152
rect 2830 1148 2834 1152
rect 2902 1158 2906 1162
rect 2982 1158 2986 1162
rect 3030 1158 3034 1162
rect 2918 1148 2922 1152
rect 2950 1148 2954 1152
rect 3014 1148 3018 1152
rect 3078 1148 3082 1152
rect 3094 1148 3098 1152
rect 3102 1148 3106 1152
rect 3118 1148 3122 1152
rect 3174 1158 3178 1162
rect 3262 1158 3266 1162
rect 3414 1158 3418 1162
rect 3158 1148 3162 1152
rect 3182 1148 3186 1152
rect 3198 1148 3202 1152
rect 3230 1148 3234 1152
rect 3246 1148 3250 1152
rect 3326 1148 3330 1152
rect 3350 1148 3354 1152
rect 3366 1148 3370 1152
rect 3382 1148 3386 1152
rect 3406 1148 3410 1152
rect 3462 1147 3466 1151
rect 3534 1148 3538 1152
rect 950 1138 954 1142
rect 974 1138 978 1142
rect 1014 1138 1018 1142
rect 1054 1138 1058 1142
rect 1094 1138 1098 1142
rect 1206 1138 1210 1142
rect 1230 1138 1234 1142
rect 1286 1138 1290 1142
rect 1342 1138 1346 1142
rect 1374 1138 1378 1142
rect 1446 1138 1450 1142
rect 1478 1138 1482 1142
rect 1526 1138 1530 1142
rect 1550 1138 1554 1142
rect 1622 1138 1626 1142
rect 1630 1138 1634 1142
rect 1662 1138 1666 1142
rect 1710 1138 1714 1142
rect 1734 1138 1738 1142
rect 1758 1138 1762 1142
rect 1806 1138 1810 1142
rect 1846 1138 1850 1142
rect 1878 1138 1882 1142
rect 1934 1138 1938 1142
rect 1958 1138 1962 1142
rect 1974 1138 1978 1142
rect 1982 1138 1986 1142
rect 2014 1138 2018 1142
rect 2070 1138 2074 1142
rect 2110 1138 2114 1142
rect 2158 1138 2162 1142
rect 2166 1138 2170 1142
rect 2182 1138 2186 1142
rect 2198 1138 2202 1142
rect 2214 1138 2218 1142
rect 2230 1138 2234 1142
rect 2246 1138 2250 1142
rect 2262 1138 2266 1142
rect 2278 1138 2282 1142
rect 2366 1138 2370 1142
rect 2406 1138 2410 1142
rect 2446 1138 2450 1142
rect 2454 1140 2458 1144
rect 2486 1138 2490 1142
rect 2502 1138 2506 1142
rect 2526 1138 2530 1142
rect 2606 1138 2610 1142
rect 2638 1138 2642 1142
rect 2702 1138 2706 1142
rect 2718 1138 2722 1142
rect 2790 1138 2794 1142
rect 2822 1138 2826 1142
rect 2878 1138 2882 1142
rect 2926 1138 2930 1142
rect 2958 1138 2962 1142
rect 2990 1138 2994 1142
rect 3006 1138 3010 1142
rect 3102 1138 3106 1142
rect 3126 1138 3130 1142
rect 3142 1138 3146 1142
rect 3150 1138 3154 1142
rect 3182 1138 3186 1142
rect 3222 1138 3226 1142
rect 3318 1138 3322 1142
rect 3350 1138 3354 1142
rect 3358 1138 3362 1142
rect 3374 1138 3378 1142
rect 3478 1138 3482 1142
rect 78 1128 82 1132
rect 254 1128 258 1132
rect 574 1128 578 1132
rect 782 1128 786 1132
rect 878 1128 882 1132
rect 926 1128 930 1132
rect 1230 1128 1234 1132
rect 1414 1128 1418 1132
rect 1718 1128 1722 1132
rect 1838 1128 1842 1132
rect 1870 1128 1874 1132
rect 1934 1128 1938 1132
rect 2006 1128 2010 1132
rect 2054 1128 2058 1132
rect 2102 1128 2106 1132
rect 2318 1128 2322 1132
rect 2350 1128 2354 1132
rect 2542 1128 2546 1132
rect 2558 1128 2562 1132
rect 2734 1128 2738 1132
rect 2766 1128 2770 1132
rect 2894 1128 2898 1132
rect 2990 1128 2994 1132
rect 3038 1128 3042 1132
rect 3078 1128 3082 1132
rect 3094 1128 3098 1132
rect 3206 1128 3210 1132
rect 3430 1128 3434 1132
rect 86 1118 90 1122
rect 118 1118 122 1122
rect 166 1118 170 1122
rect 318 1118 322 1122
rect 358 1118 362 1122
rect 430 1118 434 1122
rect 542 1118 546 1122
rect 590 1118 594 1122
rect 622 1118 626 1122
rect 734 1118 738 1122
rect 886 1118 890 1122
rect 958 1118 962 1122
rect 982 1118 986 1122
rect 1118 1118 1122 1122
rect 1406 1118 1410 1122
rect 1694 1118 1698 1122
rect 1814 1118 1818 1122
rect 2094 1118 2098 1122
rect 2358 1118 2362 1122
rect 2430 1118 2434 1122
rect 2486 1118 2490 1122
rect 2662 1118 2666 1122
rect 2814 1118 2818 1122
rect 3302 1118 3306 1122
rect 994 1103 998 1107
rect 1001 1103 1005 1107
rect 2026 1103 2030 1107
rect 2033 1103 2037 1107
rect 3042 1103 3046 1107
rect 3049 1103 3053 1107
rect 6 1088 10 1092
rect 174 1088 178 1092
rect 262 1088 266 1092
rect 398 1088 402 1092
rect 430 1088 434 1092
rect 502 1088 506 1092
rect 742 1088 746 1092
rect 830 1088 834 1092
rect 910 1088 914 1092
rect 1022 1088 1026 1092
rect 1062 1088 1066 1092
rect 1158 1088 1162 1092
rect 1222 1088 1226 1092
rect 1286 1088 1290 1092
rect 1350 1088 1354 1092
rect 1398 1088 1402 1092
rect 1502 1088 1506 1092
rect 1734 1088 1738 1092
rect 1790 1088 1794 1092
rect 1934 1088 1938 1092
rect 2006 1088 2010 1092
rect 2062 1088 2066 1092
rect 2134 1088 2138 1092
rect 2526 1088 2530 1092
rect 2694 1088 2698 1092
rect 2718 1088 2722 1092
rect 2806 1088 2810 1092
rect 2902 1088 2906 1092
rect 2982 1088 2986 1092
rect 3110 1088 3114 1092
rect 3214 1088 3218 1092
rect 3238 1088 3242 1092
rect 3294 1088 3298 1092
rect 3526 1088 3530 1092
rect 46 1078 50 1082
rect 54 1078 58 1082
rect 70 1078 74 1082
rect 110 1078 114 1082
rect 862 1078 866 1082
rect 1070 1078 1074 1082
rect 1086 1078 1090 1082
rect 1142 1078 1146 1082
rect 1174 1078 1178 1082
rect 1246 1078 1250 1082
rect 1294 1078 1298 1082
rect 1334 1078 1338 1082
rect 1454 1078 1458 1082
rect 1462 1078 1466 1082
rect 1478 1078 1482 1082
rect 1550 1078 1554 1082
rect 1614 1078 1618 1082
rect 1686 1078 1690 1082
rect 1742 1078 1746 1082
rect 1750 1078 1754 1082
rect 1798 1078 1802 1082
rect 1830 1078 1834 1082
rect 1838 1078 1842 1082
rect 1902 1078 1906 1082
rect 2054 1078 2058 1082
rect 2118 1078 2122 1082
rect 2142 1078 2146 1082
rect 2174 1078 2178 1082
rect 2246 1078 2250 1082
rect 2326 1078 2330 1082
rect 54 1068 58 1072
rect 118 1068 122 1072
rect 142 1068 146 1072
rect 198 1068 202 1072
rect 238 1068 242 1072
rect 286 1068 290 1072
rect 22 1058 26 1062
rect 86 1058 90 1062
rect 150 1058 154 1062
rect 166 1058 170 1062
rect 198 1058 202 1062
rect 206 1058 210 1062
rect 278 1058 282 1062
rect 286 1058 290 1062
rect 310 1068 314 1072
rect 342 1068 346 1072
rect 350 1068 354 1072
rect 374 1068 378 1072
rect 422 1068 426 1072
rect 454 1068 458 1072
rect 462 1068 466 1072
rect 526 1068 530 1072
rect 550 1068 554 1072
rect 566 1068 570 1072
rect 582 1068 586 1072
rect 614 1068 618 1072
rect 302 1058 306 1062
rect 374 1058 378 1062
rect 382 1058 386 1062
rect 446 1058 450 1062
rect 518 1058 522 1062
rect 574 1058 578 1062
rect 606 1058 610 1062
rect 614 1058 618 1062
rect 726 1068 730 1072
rect 750 1068 754 1072
rect 774 1068 778 1072
rect 806 1068 810 1072
rect 838 1068 842 1072
rect 878 1068 882 1072
rect 934 1068 938 1072
rect 942 1068 946 1072
rect 1038 1068 1042 1072
rect 1046 1068 1050 1072
rect 1118 1068 1122 1072
rect 1174 1068 1178 1072
rect 1222 1068 1226 1072
rect 1238 1068 1242 1072
rect 1270 1068 1274 1072
rect 1342 1068 1346 1072
rect 1374 1068 1378 1072
rect 1390 1068 1394 1072
rect 1486 1068 1490 1072
rect 1534 1068 1538 1072
rect 1550 1068 1554 1072
rect 1566 1068 1570 1072
rect 1590 1068 1594 1072
rect 1598 1068 1602 1072
rect 1654 1068 1658 1072
rect 1662 1068 1666 1072
rect 1710 1068 1714 1072
rect 1726 1068 1730 1072
rect 1782 1068 1786 1072
rect 1814 1068 1818 1072
rect 1838 1068 1842 1072
rect 1886 1068 1890 1072
rect 1910 1068 1914 1072
rect 1982 1068 1986 1072
rect 1998 1068 2002 1072
rect 2014 1068 2018 1072
rect 2030 1068 2034 1072
rect 2086 1068 2090 1072
rect 2102 1068 2106 1072
rect 2158 1068 2162 1072
rect 2206 1068 2210 1072
rect 2238 1068 2242 1072
rect 2262 1068 2266 1072
rect 2286 1068 2290 1072
rect 2398 1078 2402 1082
rect 2614 1078 2618 1082
rect 2686 1078 2690 1082
rect 2830 1078 2834 1082
rect 2910 1078 2914 1082
rect 2974 1078 2978 1082
rect 3006 1078 3010 1082
rect 3046 1078 3050 1082
rect 3086 1078 3090 1082
rect 3118 1078 3122 1082
rect 3166 1078 3170 1082
rect 3198 1078 3202 1082
rect 3286 1078 3290 1082
rect 3342 1078 3346 1082
rect 3430 1078 3434 1082
rect 2350 1068 2354 1072
rect 2430 1068 2434 1072
rect 2550 1068 2554 1072
rect 2606 1068 2610 1072
rect 2630 1068 2634 1072
rect 2638 1068 2642 1072
rect 2654 1068 2658 1072
rect 2662 1068 2666 1072
rect 2678 1068 2682 1072
rect 2702 1068 2706 1072
rect 2742 1068 2746 1072
rect 2750 1068 2754 1072
rect 2798 1068 2802 1072
rect 2846 1068 2850 1072
rect 2878 1068 2882 1072
rect 2886 1068 2890 1072
rect 2926 1068 2930 1072
rect 2990 1068 2994 1072
rect 3062 1068 3066 1072
rect 3150 1068 3154 1072
rect 3182 1068 3186 1072
rect 3254 1068 3258 1072
rect 3286 1068 3290 1072
rect 3302 1068 3306 1072
rect 3326 1068 3330 1072
rect 3350 1068 3354 1072
rect 3414 1068 3418 1072
rect 3478 1068 3482 1072
rect 646 1058 650 1062
rect 670 1058 674 1062
rect 678 1058 682 1062
rect 686 1058 690 1062
rect 710 1058 714 1062
rect 782 1058 786 1062
rect 798 1058 802 1062
rect 814 1058 818 1062
rect 886 1058 890 1062
rect 926 1058 930 1062
rect 950 1058 954 1062
rect 974 1058 978 1062
rect 982 1058 986 1062
rect 1070 1058 1074 1062
rect 1094 1058 1098 1062
rect 1126 1058 1130 1062
rect 1190 1058 1194 1062
rect 1262 1058 1266 1062
rect 1310 1058 1314 1062
rect 1350 1058 1354 1062
rect 1366 1058 1370 1062
rect 1382 1058 1386 1062
rect 1430 1058 1434 1062
rect 1462 1058 1466 1062
rect 1518 1058 1522 1062
rect 1574 1058 1578 1062
rect 1590 1058 1594 1062
rect 1630 1058 1634 1062
rect 1646 1058 1650 1062
rect 1670 1058 1674 1062
rect 1718 1058 1722 1062
rect 1766 1058 1770 1062
rect 1774 1058 1778 1062
rect 1806 1058 1810 1062
rect 1854 1058 1858 1062
rect 1886 1058 1890 1062
rect 1918 1058 1922 1062
rect 1942 1058 1946 1062
rect 1950 1058 1954 1062
rect 1974 1058 1978 1062
rect 1990 1058 1994 1062
rect 2038 1058 2042 1062
rect 2078 1058 2082 1062
rect 2094 1058 2098 1062
rect 2118 1058 2122 1062
rect 2126 1058 2130 1062
rect 2142 1058 2146 1062
rect 2150 1058 2154 1062
rect 2230 1058 2234 1062
rect 2310 1058 2314 1062
rect 2326 1058 2330 1062
rect 2358 1058 2362 1062
rect 2382 1058 2386 1062
rect 2422 1058 2426 1062
rect 2478 1058 2482 1062
rect 2494 1058 2498 1062
rect 2558 1058 2562 1062
rect 2598 1058 2602 1062
rect 2638 1058 2642 1062
rect 2646 1058 2650 1062
rect 2678 1058 2682 1062
rect 2710 1058 2714 1062
rect 2734 1058 2738 1062
rect 2806 1058 2810 1062
rect 2846 1058 2850 1062
rect 2870 1058 2874 1062
rect 2934 1058 2938 1062
rect 2950 1058 2954 1062
rect 2998 1058 3002 1062
rect 3022 1058 3026 1062
rect 3062 1058 3066 1062
rect 3094 1058 3098 1062
rect 3174 1058 3178 1062
rect 3246 1058 3250 1062
rect 3262 1058 3266 1062
rect 3310 1058 3314 1062
rect 3318 1058 3322 1062
rect 3358 1058 3362 1062
rect 3382 1058 3386 1062
rect 3398 1058 3402 1062
rect 3414 1058 3418 1062
rect 3462 1059 3466 1063
rect 6 1048 10 1052
rect 70 1048 74 1052
rect 134 1048 138 1052
rect 166 1048 170 1052
rect 174 1048 178 1052
rect 254 1048 258 1052
rect 318 1048 322 1052
rect 366 1048 370 1052
rect 398 1048 402 1052
rect 406 1048 410 1052
rect 478 1048 482 1052
rect 534 1048 538 1052
rect 590 1048 594 1052
rect 638 1048 642 1052
rect 742 1048 746 1052
rect 766 1048 770 1052
rect 798 1048 802 1052
rect 854 1048 858 1052
rect 902 1048 906 1052
rect 910 1048 914 1052
rect 966 1048 970 1052
rect 1022 1048 1026 1052
rect 1062 1048 1066 1052
rect 1150 1048 1154 1052
rect 1214 1048 1218 1052
rect 1294 1048 1298 1052
rect 1414 1048 1418 1052
rect 1502 1048 1506 1052
rect 1558 1048 1562 1052
rect 1646 1048 1650 1052
rect 1686 1048 1690 1052
rect 1694 1048 1698 1052
rect 1710 1048 1714 1052
rect 1878 1048 1882 1052
rect 2062 1048 2066 1052
rect 2182 1048 2186 1052
rect 2294 1048 2298 1052
rect 2406 1048 2410 1052
rect 2606 1048 2610 1052
rect 2718 1048 2722 1052
rect 2806 1048 2810 1052
rect 2854 1048 2858 1052
rect 2902 1048 2906 1052
rect 2934 1048 2938 1052
rect 2950 1048 2954 1052
rect 3126 1048 3130 1052
rect 3158 1048 3162 1052
rect 3206 1048 3210 1052
rect 3230 1048 3234 1052
rect 3278 1048 3282 1052
rect 3342 1048 3346 1052
rect 3374 1048 3378 1052
rect 126 1038 130 1042
rect 342 1038 346 1042
rect 1334 1038 1338 1042
rect 2174 1038 2178 1042
rect 2766 1038 2770 1042
rect 3174 1038 3178 1042
rect 3558 1038 3562 1042
rect 1262 1028 1266 1032
rect 3142 1028 3146 1032
rect 606 1018 610 1022
rect 630 1018 634 1022
rect 702 1018 706 1022
rect 758 1018 762 1022
rect 870 1018 874 1022
rect 886 1018 890 1022
rect 950 1018 954 1022
rect 1006 1018 1010 1022
rect 1134 1018 1138 1022
rect 1182 1018 1186 1022
rect 1278 1018 1282 1022
rect 1758 1018 1762 1022
rect 1886 1018 1890 1022
rect 2198 1018 2202 1022
rect 2334 1018 2338 1022
rect 2358 1018 2362 1022
rect 2422 1018 2426 1022
rect 2558 1018 2562 1022
rect 2918 1018 2922 1022
rect 482 1003 486 1007
rect 489 1003 493 1007
rect 1514 1003 1518 1007
rect 1521 1003 1525 1007
rect 2538 1003 2542 1007
rect 2545 1003 2549 1007
rect 30 988 34 992
rect 126 988 130 992
rect 302 988 306 992
rect 446 988 450 992
rect 470 988 474 992
rect 510 988 514 992
rect 590 988 594 992
rect 750 988 754 992
rect 774 988 778 992
rect 958 988 962 992
rect 1350 988 1354 992
rect 1438 988 1442 992
rect 1566 988 1570 992
rect 1598 988 1602 992
rect 1670 988 1674 992
rect 1734 988 1738 992
rect 1782 988 1786 992
rect 1878 988 1882 992
rect 1942 988 1946 992
rect 2062 988 2066 992
rect 2094 988 2098 992
rect 2246 988 2250 992
rect 2302 988 2306 992
rect 2438 988 2442 992
rect 2486 988 2490 992
rect 2590 988 2594 992
rect 2718 988 2722 992
rect 2830 988 2834 992
rect 2846 988 2850 992
rect 3206 988 3210 992
rect 3406 988 3410 992
rect 3526 988 3530 992
rect 3558 988 3562 992
rect 1318 978 1322 982
rect 3422 978 3426 982
rect 190 968 194 972
rect 230 968 234 972
rect 1646 968 1650 972
rect 3190 968 3194 972
rect 3342 968 3346 972
rect 3398 968 3402 972
rect 6 958 10 962
rect 86 958 90 962
rect 102 958 106 962
rect 110 958 114 962
rect 150 958 154 962
rect 158 958 162 962
rect 206 958 210 962
rect 270 958 274 962
rect 310 958 314 962
rect 358 958 362 962
rect 382 958 386 962
rect 414 958 418 962
rect 542 958 546 962
rect 550 958 554 962
rect 630 958 634 962
rect 694 958 698 962
rect 734 958 738 962
rect 806 958 810 962
rect 878 958 882 962
rect 70 948 74 952
rect 86 948 90 952
rect 182 948 186 952
rect 254 948 258 952
rect 270 948 274 952
rect 326 948 330 952
rect 398 948 402 952
rect 422 948 426 952
rect 430 948 434 952
rect 454 948 458 952
rect 526 948 530 952
rect 566 948 570 952
rect 622 948 626 952
rect 646 948 650 952
rect 702 948 706 952
rect 726 948 730 952
rect 750 948 754 952
rect 814 948 818 952
rect 822 948 826 952
rect 846 948 850 952
rect 942 958 946 962
rect 974 958 978 962
rect 902 948 906 952
rect 926 948 930 952
rect 958 948 962 952
rect 990 948 994 952
rect 1030 958 1034 962
rect 1102 958 1106 962
rect 1134 958 1138 962
rect 1334 958 1338 962
rect 1046 948 1050 952
rect 1062 948 1066 952
rect 1118 948 1122 952
rect 1150 948 1154 952
rect 1182 948 1186 952
rect 1214 948 1218 952
rect 1238 948 1242 952
rect 1246 948 1250 952
rect 1262 948 1266 952
rect 1270 948 1274 952
rect 1278 948 1282 952
rect 1286 948 1290 952
rect 1302 948 1306 952
rect 1318 948 1322 952
rect 1350 948 1354 952
rect 1366 948 1370 952
rect 1414 948 1418 952
rect 1430 948 1434 952
rect 1446 948 1450 952
rect 1470 948 1474 952
rect 1494 958 1498 962
rect 1614 958 1618 962
rect 1894 958 1898 962
rect 2006 958 2010 962
rect 2110 958 2114 962
rect 2454 958 2458 962
rect 2862 958 2866 962
rect 1510 948 1514 952
rect 1542 948 1546 952
rect 1550 948 1554 952
rect 1582 948 1586 952
rect 1598 948 1602 952
rect 1686 948 1690 952
rect 1718 948 1722 952
rect 1750 948 1754 952
rect 1766 948 1770 952
rect 1790 948 1794 952
rect 1798 948 1802 952
rect 1830 948 1834 952
rect 1870 948 1874 952
rect 1918 948 1922 952
rect 1966 948 1970 952
rect 1998 948 2002 952
rect 2054 948 2058 952
rect 2070 948 2074 952
rect 2094 948 2098 952
rect 2118 948 2122 952
rect 2142 948 2146 952
rect 2166 948 2170 952
rect 2182 948 2186 952
rect 2230 948 2234 952
rect 2278 948 2282 952
rect 2334 948 2338 952
rect 2382 948 2386 952
rect 2534 948 2538 952
rect 2574 948 2578 952
rect 2606 948 2610 952
rect 2638 948 2642 952
rect 2718 948 2722 952
rect 2734 948 2738 952
rect 2774 948 2778 952
rect 2782 948 2786 952
rect 2806 948 2810 952
rect 2846 948 2850 952
rect 2894 948 2898 952
rect 2918 958 2922 962
rect 2934 958 2938 962
rect 2966 958 2970 962
rect 3158 958 3162 962
rect 2942 948 2946 952
rect 2982 948 2986 952
rect 3054 948 3058 952
rect 3078 948 3082 952
rect 3094 948 3098 952
rect 3134 948 3138 952
rect 3174 948 3178 952
rect 3190 948 3194 952
rect 3214 948 3218 952
rect 3246 948 3250 952
rect 22 938 26 942
rect 94 938 98 942
rect 134 938 138 942
rect 166 938 170 942
rect 182 938 186 942
rect 222 938 226 942
rect 246 938 250 942
rect 326 938 330 942
rect 334 938 338 942
rect 350 938 354 942
rect 366 938 370 942
rect 390 938 394 942
rect 406 938 410 942
rect 518 938 522 942
rect 558 938 562 942
rect 574 938 578 942
rect 678 938 682 942
rect 758 938 762 942
rect 790 938 794 942
rect 862 938 866 942
rect 878 938 882 942
rect 910 938 914 942
rect 918 938 922 942
rect 950 938 954 942
rect 982 938 986 942
rect 1054 938 1058 942
rect 1086 938 1090 942
rect 1110 938 1114 942
rect 1126 938 1130 942
rect 1174 938 1178 942
rect 1254 938 1258 942
rect 1286 938 1290 942
rect 1294 938 1298 942
rect 1326 938 1330 942
rect 1358 938 1362 942
rect 1382 938 1386 942
rect 1422 938 1426 942
rect 1454 938 1458 942
rect 1462 938 1466 942
rect 1518 938 1522 942
rect 1582 938 1586 942
rect 1622 938 1626 942
rect 1694 938 1698 942
rect 1806 938 1810 942
rect 1854 940 1858 944
rect 1862 938 1866 942
rect 1910 938 1914 942
rect 1942 938 1946 942
rect 1958 938 1962 942
rect 2022 938 2026 942
rect 2046 938 2050 942
rect 2078 938 2082 942
rect 2086 938 2090 942
rect 2174 938 2178 942
rect 2342 938 2346 942
rect 2366 940 2370 944
rect 2374 938 2378 942
rect 2406 938 2410 942
rect 2446 938 2450 942
rect 2470 938 2474 942
rect 2478 938 2482 942
rect 2654 938 2658 942
rect 2662 938 2666 942
rect 2710 938 2714 942
rect 2742 938 2746 942
rect 2774 938 2778 942
rect 2910 938 2914 942
rect 2934 938 2938 942
rect 2974 938 2978 942
rect 2990 938 2994 942
rect 2998 938 3002 942
rect 3046 938 3050 942
rect 3086 938 3090 942
rect 3110 938 3114 942
rect 3142 938 3146 942
rect 3166 938 3170 942
rect 3278 947 3282 951
rect 3310 948 3314 952
rect 3350 948 3354 952
rect 3366 948 3370 952
rect 3382 948 3386 952
rect 3406 948 3410 952
rect 3462 947 3466 951
rect 3534 948 3538 952
rect 3198 938 3202 942
rect 3222 938 3226 942
rect 3230 938 3234 942
rect 3238 938 3242 942
rect 3350 938 3354 942
rect 3374 938 3378 942
rect 3446 938 3450 942
rect 38 928 42 932
rect 46 928 50 932
rect 118 928 122 932
rect 190 928 194 932
rect 230 928 234 932
rect 286 928 290 932
rect 294 928 298 932
rect 478 928 482 932
rect 502 928 506 932
rect 542 928 546 932
rect 582 928 586 932
rect 606 928 610 932
rect 670 928 674 932
rect 782 928 786 932
rect 1078 928 1082 932
rect 1198 928 1202 932
rect 1382 928 1386 932
rect 1886 928 1890 932
rect 1934 928 1938 932
rect 1942 928 1946 932
rect 2182 928 2186 932
rect 2198 928 2202 932
rect 2238 928 2242 932
rect 2734 928 2738 932
rect 2798 928 2802 932
rect 2830 928 2834 932
rect 2870 928 2874 932
rect 2958 928 2962 932
rect 3070 928 3074 932
rect 3102 928 3106 932
rect 3158 928 3162 932
rect 3430 928 3434 932
rect 3510 928 3514 932
rect 14 918 18 922
rect 150 918 154 922
rect 214 918 218 922
rect 270 918 274 922
rect 318 918 322 922
rect 382 918 386 922
rect 630 918 634 922
rect 694 918 698 922
rect 806 918 810 922
rect 838 918 842 922
rect 942 918 946 922
rect 1022 918 1026 922
rect 1070 918 1074 922
rect 1102 918 1106 922
rect 1190 918 1194 922
rect 1230 918 1234 922
rect 1374 918 1378 922
rect 1398 918 1402 922
rect 1486 918 1490 922
rect 1670 918 1674 922
rect 1838 918 1842 922
rect 1902 918 1906 922
rect 1982 918 1986 922
rect 2014 918 2018 922
rect 2150 918 2154 922
rect 2262 918 2266 922
rect 2302 918 2306 922
rect 2318 918 2322 922
rect 2350 918 2354 922
rect 2462 918 2466 922
rect 2502 918 2506 922
rect 2550 918 2554 922
rect 2622 918 2626 922
rect 2694 918 2698 922
rect 2950 918 2954 922
rect 994 903 998 907
rect 1001 903 1005 907
rect 2026 903 2030 907
rect 2033 903 2037 907
rect 3042 903 3046 907
rect 3049 903 3053 907
rect 38 888 42 892
rect 142 888 146 892
rect 310 888 314 892
rect 342 888 346 892
rect 374 888 378 892
rect 414 888 418 892
rect 478 888 482 892
rect 534 888 538 892
rect 550 888 554 892
rect 654 888 658 892
rect 734 888 738 892
rect 886 888 890 892
rect 942 888 946 892
rect 974 888 978 892
rect 1094 888 1098 892
rect 1134 888 1138 892
rect 1166 888 1170 892
rect 1214 888 1218 892
rect 1366 888 1370 892
rect 1414 888 1418 892
rect 1670 888 1674 892
rect 1686 888 1690 892
rect 1782 888 1786 892
rect 2190 888 2194 892
rect 2270 888 2274 892
rect 2454 888 2458 892
rect 2710 888 2714 892
rect 2742 888 2746 892
rect 2806 888 2810 892
rect 2846 888 2850 892
rect 2966 888 2970 892
rect 3102 888 3106 892
rect 3134 888 3138 892
rect 3166 888 3170 892
rect 3246 888 3250 892
rect 3254 888 3258 892
rect 3302 888 3306 892
rect 3358 888 3362 892
rect 3406 888 3410 892
rect 3438 888 3442 892
rect 182 878 186 882
rect 286 878 290 882
rect 462 878 466 882
rect 478 878 482 882
rect 622 878 626 882
rect 1054 878 1058 882
rect 1158 878 1162 882
rect 1246 878 1250 882
rect 1270 878 1274 882
rect 1422 878 1426 882
rect 1518 878 1522 882
rect 1534 878 1538 882
rect 6 868 10 872
rect 62 868 66 872
rect 86 868 90 872
rect 94 868 98 872
rect 110 868 114 872
rect 198 868 202 872
rect 214 868 218 872
rect 230 868 234 872
rect 246 868 250 872
rect 254 868 258 872
rect 334 868 338 872
rect 366 868 370 872
rect 398 868 402 872
rect 422 868 426 872
rect 438 868 442 872
rect 462 868 466 872
rect 518 868 522 872
rect 542 868 546 872
rect 574 868 578 872
rect 606 868 610 872
rect 630 868 634 872
rect 686 868 690 872
rect 702 868 706 872
rect 718 868 722 872
rect 750 868 754 872
rect 766 868 770 872
rect 798 868 802 872
rect 806 868 810 872
rect 910 868 914 872
rect 990 868 994 872
rect 1014 868 1018 872
rect 1038 868 1042 872
rect 1062 868 1066 872
rect 1118 868 1122 872
rect 1142 868 1146 872
rect 1182 868 1186 872
rect 1190 868 1194 872
rect 1230 868 1234 872
rect 1254 868 1258 872
rect 1302 868 1306 872
rect 38 858 42 862
rect 62 858 66 862
rect 158 858 162 862
rect 206 858 210 862
rect 238 858 242 862
rect 302 858 306 862
rect 326 858 330 862
rect 358 858 362 862
rect 390 858 394 862
rect 446 858 450 862
rect 510 858 514 862
rect 566 858 570 862
rect 598 858 602 862
rect 622 858 626 862
rect 686 858 690 862
rect 718 858 722 862
rect 790 858 794 862
rect 814 858 818 862
rect 838 858 842 862
rect 846 858 850 862
rect 870 858 874 862
rect 902 858 906 862
rect 926 858 930 862
rect 950 858 954 862
rect 966 858 970 862
rect 1030 858 1034 862
rect 1070 858 1074 862
rect 1110 858 1114 862
rect 1182 858 1186 862
rect 1222 858 1226 862
rect 1254 858 1258 862
rect 1294 858 1298 862
rect 1302 858 1306 862
rect 1398 868 1402 872
rect 1438 868 1442 872
rect 1454 868 1458 872
rect 1470 868 1474 872
rect 1486 868 1490 872
rect 1542 868 1546 872
rect 1590 868 1594 872
rect 2294 878 2298 882
rect 2310 878 2314 882
rect 2462 878 2466 882
rect 2526 878 2530 882
rect 2734 878 2738 882
rect 1622 868 1626 872
rect 1646 868 1650 872
rect 1694 868 1698 872
rect 1702 868 1706 872
rect 1758 868 1762 872
rect 1798 868 1802 872
rect 1318 858 1322 862
rect 1350 858 1354 862
rect 1390 858 1394 862
rect 1406 858 1410 862
rect 1446 858 1450 862
rect 1478 858 1482 862
rect 1494 858 1498 862
rect 1582 858 1586 862
rect 1614 858 1618 862
rect 1638 858 1642 862
rect 1726 858 1730 862
rect 1766 858 1770 862
rect 1806 858 1810 862
rect 1822 858 1826 862
rect 1846 858 1850 862
rect 1886 868 1890 872
rect 1918 868 1922 872
rect 1950 868 1954 872
rect 1958 868 1962 872
rect 1974 868 1978 872
rect 2006 868 2010 872
rect 2054 868 2058 872
rect 2062 868 2066 872
rect 2118 868 2122 872
rect 2134 868 2138 872
rect 2150 868 2154 872
rect 2166 868 2170 872
rect 2174 866 2178 870
rect 2198 868 2202 872
rect 2230 868 2234 872
rect 2278 868 2282 872
rect 2318 868 2322 872
rect 2350 868 2354 872
rect 2374 868 2378 872
rect 2390 868 2394 872
rect 2430 868 2434 872
rect 2446 868 2450 872
rect 2510 868 2514 872
rect 2598 868 2602 872
rect 2670 868 2674 872
rect 2814 878 2818 882
rect 2830 878 2834 882
rect 3070 878 3074 882
rect 3126 878 3130 882
rect 3158 878 3162 882
rect 3182 878 3186 882
rect 3214 878 3218 882
rect 2750 868 2754 872
rect 2766 868 2770 872
rect 2774 868 2778 872
rect 2790 868 2794 872
rect 2854 868 2858 872
rect 2926 868 2930 872
rect 2942 868 2946 872
rect 2950 868 2954 872
rect 2974 868 2978 872
rect 3038 868 3042 872
rect 3078 868 3082 872
rect 3214 868 3218 872
rect 3278 868 3282 872
rect 3286 868 3290 872
rect 3334 868 3338 872
rect 3342 868 3346 872
rect 3390 868 3394 872
rect 3398 868 3402 872
rect 3494 868 3498 872
rect 3518 868 3522 872
rect 1878 858 1882 862
rect 1894 858 1898 862
rect 1950 858 1954 862
rect 1998 858 2002 862
rect 2038 858 2042 862
rect 2054 858 2058 862
rect 2062 858 2066 862
rect 2086 858 2090 862
rect 2110 858 2114 862
rect 2126 858 2130 862
rect 2158 858 2162 862
rect 2206 858 2210 862
rect 2222 858 2226 862
rect 2286 858 2290 862
rect 2294 858 2298 862
rect 2326 858 2330 862
rect 2358 858 2362 862
rect 2382 858 2386 862
rect 2438 858 2442 862
rect 2486 858 2490 862
rect 2502 858 2506 862
rect 2518 858 2522 862
rect 2574 858 2578 862
rect 2670 858 2674 862
rect 2750 858 2754 862
rect 2830 858 2834 862
rect 2870 858 2874 862
rect 2902 858 2906 862
rect 2982 858 2986 862
rect 3022 858 3026 862
rect 3030 858 3034 862
rect 3046 858 3050 862
rect 3086 858 3090 862
rect 3110 858 3114 862
rect 3174 858 3178 862
rect 3230 858 3234 862
rect 3286 858 3290 862
rect 3422 858 3426 862
rect 3502 858 3506 862
rect 3526 858 3530 862
rect 38 848 42 852
rect 70 848 74 852
rect 86 848 90 852
rect 118 848 122 852
rect 142 848 146 852
rect 190 848 194 852
rect 222 848 226 852
rect 270 848 274 852
rect 310 848 314 852
rect 342 848 346 852
rect 374 848 378 852
rect 406 848 410 852
rect 430 848 434 852
rect 494 848 498 852
rect 526 848 530 852
rect 550 848 554 852
rect 582 848 586 852
rect 654 848 658 852
rect 662 848 666 852
rect 694 848 698 852
rect 726 848 730 852
rect 750 848 754 852
rect 774 848 778 852
rect 830 848 834 852
rect 886 848 890 852
rect 966 848 970 852
rect 990 848 994 852
rect 1054 848 1058 852
rect 1086 848 1090 852
rect 1094 848 1098 852
rect 1126 848 1130 852
rect 1158 848 1162 852
rect 1214 848 1218 852
rect 1278 848 1282 852
rect 1334 848 1338 852
rect 1366 848 1370 852
rect 1374 848 1378 852
rect 1390 848 1394 852
rect 1430 848 1434 852
rect 1462 848 1466 852
rect 1566 848 1570 852
rect 1582 848 1586 852
rect 1670 848 1674 852
rect 1678 848 1682 852
rect 1726 848 1730 852
rect 1830 848 1834 852
rect 1926 848 1930 852
rect 1974 848 1978 852
rect 1982 848 1986 852
rect 2014 848 2018 852
rect 2086 848 2090 852
rect 2110 848 2114 852
rect 2222 848 2226 852
rect 2254 848 2258 852
rect 2342 848 2346 852
rect 2414 848 2418 852
rect 2494 848 2498 852
rect 2694 848 2698 852
rect 2710 848 2714 852
rect 2806 848 2810 852
rect 2838 848 2842 852
rect 2886 848 2890 852
rect 2918 848 2922 852
rect 2926 848 2930 852
rect 2966 848 2970 852
rect 2998 848 3002 852
rect 3134 848 3138 852
rect 3254 848 3258 852
rect 54 838 58 842
rect 94 838 98 842
rect 118 838 122 842
rect 254 838 258 842
rect 1158 838 1162 842
rect 1558 838 1562 842
rect 2326 838 2330 842
rect 2478 838 2482 842
rect 3022 838 3026 842
rect 3558 838 3562 842
rect 598 828 602 832
rect 614 828 618 832
rect 758 828 762 832
rect 1262 828 1266 832
rect 1638 828 1642 832
rect 2590 828 2594 832
rect 678 818 682 822
rect 790 818 794 822
rect 814 818 818 822
rect 862 818 866 822
rect 998 818 1002 822
rect 1070 818 1074 822
rect 1294 818 1298 822
rect 1502 818 1506 822
rect 1710 818 1714 822
rect 1750 818 1754 822
rect 1846 818 1850 822
rect 1910 818 1914 822
rect 1942 818 1946 822
rect 1998 818 2002 822
rect 2150 818 2154 822
rect 2206 818 2210 822
rect 2406 818 2410 822
rect 2486 818 2490 822
rect 2558 818 2562 822
rect 2614 818 2618 822
rect 2782 818 2786 822
rect 3438 818 3442 822
rect 482 803 486 807
rect 489 803 493 807
rect 1514 803 1518 807
rect 1521 803 1525 807
rect 2538 803 2542 807
rect 2545 803 2549 807
rect 54 788 58 792
rect 126 788 130 792
rect 150 788 154 792
rect 174 788 178 792
rect 198 788 202 792
rect 214 788 218 792
rect 238 788 242 792
rect 398 788 402 792
rect 422 788 426 792
rect 598 788 602 792
rect 726 788 730 792
rect 742 788 746 792
rect 806 788 810 792
rect 846 788 850 792
rect 1086 788 1090 792
rect 1166 788 1170 792
rect 1310 788 1314 792
rect 1366 788 1370 792
rect 1406 788 1410 792
rect 1454 788 1458 792
rect 1518 788 1522 792
rect 1790 788 1794 792
rect 1838 788 1842 792
rect 2678 788 2682 792
rect 3062 788 3066 792
rect 3126 788 3130 792
rect 3422 788 3426 792
rect 3470 788 3474 792
rect 3494 788 3498 792
rect 3550 788 3554 792
rect 582 778 586 782
rect 2638 778 2642 782
rect 2950 778 2954 782
rect 3102 778 3106 782
rect 3518 778 3522 782
rect 870 768 874 772
rect 1246 768 1250 772
rect 1398 768 1402 772
rect 1478 768 1482 772
rect 1534 768 1538 772
rect 1566 768 1570 772
rect 2598 768 2602 772
rect 2790 768 2794 772
rect 3094 768 3098 772
rect 3182 768 3186 772
rect 94 758 98 762
rect 158 758 162 762
rect 222 758 226 762
rect 262 758 266 762
rect 270 758 274 762
rect 302 758 306 762
rect 318 758 322 762
rect 350 758 354 762
rect 374 758 378 762
rect 30 748 34 752
rect 78 748 82 752
rect 174 748 178 752
rect 286 748 290 752
rect 318 748 322 752
rect 398 748 402 752
rect 446 758 450 762
rect 502 758 506 762
rect 590 758 594 762
rect 638 758 642 762
rect 526 748 530 752
rect 558 748 562 752
rect 566 748 570 752
rect 622 748 626 752
rect 718 758 722 762
rect 702 748 706 752
rect 742 748 746 752
rect 766 758 770 762
rect 814 758 818 762
rect 886 758 890 762
rect 918 758 922 762
rect 926 758 930 762
rect 950 758 954 762
rect 998 758 1002 762
rect 782 748 786 752
rect 822 748 826 752
rect 830 748 834 752
rect 854 748 858 752
rect 886 748 890 752
rect 902 748 906 752
rect 926 748 930 752
rect 982 748 986 752
rect 1078 758 1082 762
rect 1118 758 1122 762
rect 1150 758 1154 762
rect 1222 758 1226 762
rect 1230 758 1234 762
rect 1286 758 1290 762
rect 1414 758 1418 762
rect 1062 748 1066 752
rect 1126 748 1130 752
rect 1150 748 1154 752
rect 1166 748 1170 752
rect 1206 748 1210 752
rect 1214 748 1218 752
rect 1246 748 1250 752
rect 1270 748 1274 752
rect 1278 748 1282 752
rect 1294 748 1298 752
rect 1302 748 1306 752
rect 1334 748 1338 752
rect 1342 748 1346 752
rect 1350 748 1354 752
rect 1374 748 1378 752
rect 1406 748 1410 752
rect 1422 748 1426 752
rect 1486 758 1490 762
rect 1606 758 1610 762
rect 1630 758 1634 762
rect 1638 758 1642 762
rect 1814 758 1818 762
rect 1854 758 1858 762
rect 1910 758 1914 762
rect 1486 748 1490 752
rect 1550 748 1554 752
rect 1590 748 1594 752
rect 1614 748 1618 752
rect 1686 748 1690 752
rect 1694 748 1698 752
rect 1742 748 1746 752
rect 1766 748 1770 752
rect 1774 748 1778 752
rect 1838 748 1842 752
rect 1862 748 1866 752
rect 2006 758 2010 762
rect 2014 758 2018 762
rect 2094 758 2098 762
rect 2142 758 2146 762
rect 2158 758 2162 762
rect 2422 758 2426 762
rect 2454 758 2458 762
rect 2654 758 2658 762
rect 2822 758 2826 762
rect 1934 748 1938 752
rect 1990 748 1994 752
rect 2078 748 2082 752
rect 2118 748 2122 752
rect 2134 748 2138 752
rect 2166 748 2170 752
rect 2198 748 2202 752
rect 2222 748 2226 752
rect 2246 748 2250 752
rect 2254 748 2258 752
rect 2286 748 2290 752
rect 2342 747 2346 751
rect 2374 748 2378 752
rect 2414 748 2418 752
rect 2462 748 2466 752
rect 2494 748 2498 752
rect 2534 747 2538 751
rect 2606 748 2610 752
rect 2630 748 2634 752
rect 2734 748 2738 752
rect 2742 748 2746 752
rect 2798 748 2802 752
rect 2806 748 2810 752
rect 2846 758 2850 762
rect 3078 758 3082 762
rect 3110 758 3114 762
rect 3118 758 3122 762
rect 3166 758 3170 762
rect 2854 748 2858 752
rect 2886 747 2890 751
rect 2958 748 2962 752
rect 2982 748 2986 752
rect 3030 748 3034 752
rect 3054 748 3058 752
rect 3102 748 3106 752
rect 3142 748 3146 752
rect 3182 748 3186 752
rect 3214 748 3218 752
rect 3230 748 3234 752
rect 3262 747 3266 751
rect 3294 748 3298 752
rect 3358 747 3362 751
rect 3390 748 3394 752
rect 3430 748 3434 752
rect 3454 748 3458 752
rect 3478 748 3482 752
rect 3502 748 3506 752
rect 3526 748 3530 752
rect 38 738 42 742
rect 70 738 74 742
rect 86 738 90 742
rect 134 738 138 742
rect 182 738 186 742
rect 206 738 210 742
rect 246 738 250 742
rect 262 738 266 742
rect 294 738 298 742
rect 326 738 330 742
rect 334 738 338 742
rect 358 738 362 742
rect 406 738 410 742
rect 414 738 418 742
rect 462 738 466 742
rect 518 738 522 742
rect 574 738 578 742
rect 614 738 618 742
rect 630 738 634 742
rect 662 738 666 742
rect 678 738 682 742
rect 694 738 698 742
rect 734 738 738 742
rect 790 738 794 742
rect 798 738 802 742
rect 870 738 874 742
rect 894 738 898 742
rect 942 738 946 742
rect 966 738 970 742
rect 974 738 978 742
rect 1038 738 1042 742
rect 1054 738 1058 742
rect 1070 738 1074 742
rect 1094 738 1098 742
rect 1102 738 1106 742
rect 1254 738 1258 742
rect 1262 738 1266 742
rect 1326 738 1330 742
rect 1462 738 1466 742
rect 1574 738 1578 742
rect 1614 738 1618 742
rect 1654 738 1658 742
rect 1670 738 1674 742
rect 1734 738 1738 742
rect 1822 738 1826 742
rect 1830 738 1834 742
rect 1878 738 1882 742
rect 1886 738 1890 742
rect 1926 738 1930 742
rect 1942 738 1946 742
rect 1958 738 1962 742
rect 1982 738 1986 742
rect 2030 738 2034 742
rect 2070 738 2074 742
rect 2126 738 2130 742
rect 2134 738 2138 742
rect 2174 738 2178 742
rect 2230 738 2234 742
rect 2262 738 2266 742
rect 2278 738 2282 742
rect 2294 738 2298 742
rect 2310 738 2314 742
rect 2438 738 2442 742
rect 2454 738 2458 742
rect 2470 738 2474 742
rect 2542 738 2546 742
rect 2550 738 2554 742
rect 2606 738 2610 742
rect 2630 738 2634 742
rect 2662 738 2666 742
rect 2710 738 2714 742
rect 2750 738 2754 742
rect 2774 738 2778 742
rect 2798 738 2802 742
rect 2854 738 2858 742
rect 2870 738 2874 742
rect 2974 738 2978 742
rect 3022 738 3026 742
rect 3054 738 3058 742
rect 3190 738 3194 742
rect 3230 738 3234 742
rect 3446 738 3450 742
rect 38 728 42 732
rect 62 728 66 732
rect 142 728 146 732
rect 190 728 194 732
rect 230 728 234 732
rect 470 728 474 732
rect 606 728 610 732
rect 702 728 706 732
rect 718 728 722 732
rect 1142 728 1146 732
rect 1182 728 1186 732
rect 1438 728 1442 732
rect 1502 728 1506 732
rect 1518 728 1522 732
rect 1662 728 1666 732
rect 1710 728 1714 732
rect 1750 728 1754 732
rect 1950 728 1954 732
rect 2006 728 2010 732
rect 2054 728 2058 732
rect 2094 728 2098 732
rect 2214 728 2218 732
rect 2246 728 2250 732
rect 2278 728 2282 732
rect 2310 728 2314 732
rect 2430 728 2434 732
rect 2486 728 2490 732
rect 2622 728 2626 732
rect 2718 728 2722 732
rect 2766 728 2770 732
rect 2774 728 2778 732
rect 2966 728 2970 732
rect 3006 728 3010 732
rect 3158 728 3162 732
rect 3198 728 3202 732
rect 14 718 18 722
rect 342 718 346 722
rect 486 718 490 722
rect 510 718 514 722
rect 542 718 546 722
rect 934 718 938 722
rect 958 718 962 722
rect 1006 718 1010 722
rect 1110 718 1114 722
rect 1470 718 1474 722
rect 1622 718 1626 722
rect 1646 718 1650 722
rect 1726 718 1730 722
rect 1758 718 1762 722
rect 1974 718 1978 722
rect 2014 718 2018 722
rect 2062 718 2066 722
rect 2102 718 2106 722
rect 2182 718 2186 722
rect 2406 718 2410 722
rect 2726 718 2730 722
rect 2998 718 3002 722
rect 3014 718 3018 722
rect 3206 718 3210 722
rect 3326 718 3330 722
rect 3422 718 3426 722
rect 994 703 998 707
rect 1001 703 1005 707
rect 2026 703 2030 707
rect 2033 703 2037 707
rect 3042 703 3046 707
rect 3049 703 3053 707
rect 118 688 122 692
rect 158 688 162 692
rect 190 688 194 692
rect 230 688 234 692
rect 254 688 258 692
rect 318 688 322 692
rect 398 688 402 692
rect 430 688 434 692
rect 454 688 458 692
rect 462 688 466 692
rect 494 688 498 692
rect 534 688 538 692
rect 582 688 586 692
rect 622 688 626 692
rect 654 688 658 692
rect 958 688 962 692
rect 1030 688 1034 692
rect 1046 688 1050 692
rect 1246 688 1250 692
rect 1270 688 1274 692
rect 1470 688 1474 692
rect 1566 688 1570 692
rect 1590 688 1594 692
rect 1718 688 1722 692
rect 1814 688 1818 692
rect 1862 688 1866 692
rect 1942 688 1946 692
rect 2110 688 2114 692
rect 2158 688 2162 692
rect 2318 688 2322 692
rect 2334 688 2338 692
rect 2638 688 2642 692
rect 2806 688 2810 692
rect 2846 688 2850 692
rect 2958 688 2962 692
rect 3142 688 3146 692
rect 3174 688 3178 692
rect 3198 688 3202 692
rect 3318 688 3322 692
rect 3518 688 3522 692
rect 390 678 394 682
rect 726 678 730 682
rect 830 678 834 682
rect 862 678 866 682
rect 918 678 922 682
rect 1038 678 1042 682
rect 1078 678 1082 682
rect 1262 678 1266 682
rect 1358 678 1362 682
rect 1518 678 1522 682
rect 1550 678 1554 682
rect 1574 678 1578 682
rect 1614 678 1618 682
rect 1726 678 1730 682
rect 1766 678 1770 682
rect 1822 678 1826 682
rect 1846 678 1850 682
rect 1870 678 1874 682
rect 1910 678 1914 682
rect 2166 678 2170 682
rect 14 668 18 672
rect 38 668 42 672
rect 70 668 74 672
rect 86 668 90 672
rect 94 668 98 672
rect 142 668 146 672
rect 150 668 154 672
rect 198 668 202 672
rect 294 668 298 672
rect 358 668 362 672
rect 366 668 370 672
rect 406 668 410 672
rect 438 668 442 672
rect 478 668 482 672
rect 526 668 530 672
rect 558 668 562 672
rect 566 668 570 672
rect 614 668 618 672
rect 646 668 650 672
rect 670 668 674 672
rect 758 668 762 672
rect 766 668 770 672
rect 838 668 842 672
rect 894 668 898 672
rect 918 668 922 672
rect 950 668 954 672
rect 982 668 986 672
rect 1006 668 1010 672
rect 1070 668 1074 672
rect 1086 668 1090 672
rect 1118 668 1122 672
rect 1134 668 1138 672
rect 1142 668 1146 672
rect 1198 668 1202 672
rect 1206 668 1210 672
rect 1254 668 1258 672
rect 1294 668 1298 672
rect 1310 668 1314 672
rect 1334 668 1338 672
rect 1390 668 1394 672
rect 1422 668 1426 672
rect 1430 668 1434 672
rect 1478 668 1482 672
rect 1494 668 1498 672
rect 1670 668 1674 672
rect 1710 668 1714 672
rect 1742 668 1746 672
rect 1782 668 1786 672
rect 1854 668 1858 672
rect 1902 668 1906 672
rect 1950 668 1954 672
rect 1958 668 1962 672
rect 2006 668 2010 672
rect 2030 668 2034 672
rect 2078 668 2082 672
rect 2086 668 2090 672
rect 2182 668 2186 672
rect 2206 678 2210 682
rect 2342 678 2346 682
rect 2350 678 2354 682
rect 2430 678 2434 682
rect 2510 678 2514 682
rect 2630 678 2634 682
rect 2654 678 2658 682
rect 2662 678 2666 682
rect 2710 678 2714 682
rect 2742 678 2746 682
rect 2926 678 2930 682
rect 3102 678 3106 682
rect 3150 678 3154 682
rect 3334 678 3338 682
rect 3422 678 3426 682
rect 2374 668 2378 672
rect 2414 668 2418 672
rect 2438 668 2442 672
rect 2494 668 2498 672
rect 2542 668 2546 672
rect 2670 668 2674 672
rect 2694 668 2698 672
rect 2814 668 2818 672
rect 2862 668 2866 672
rect 2894 668 2898 672
rect 2942 668 2946 672
rect 2982 668 2986 672
rect 2998 668 3002 672
rect 3006 668 3010 672
rect 3014 668 3018 672
rect 3086 668 3090 672
rect 3110 668 3114 672
rect 3166 668 3170 672
rect 3182 668 3186 672
rect 3334 668 3338 672
rect 3350 668 3354 672
rect 3366 668 3370 672
rect 3422 668 3426 672
rect 3438 668 3442 672
rect 30 658 34 662
rect 78 658 82 662
rect 134 658 138 662
rect 174 658 178 662
rect 214 658 218 662
rect 238 658 242 662
rect 294 658 298 662
rect 302 658 306 662
rect 334 658 338 662
rect 414 658 418 662
rect 518 658 522 662
rect 550 658 554 662
rect 606 658 610 662
rect 638 658 642 662
rect 678 658 682 662
rect 702 658 706 662
rect 750 658 754 662
rect 806 658 810 662
rect 846 658 850 662
rect 886 658 890 662
rect 894 658 898 662
rect 918 658 922 662
rect 958 658 962 662
rect 982 658 986 662
rect 1014 658 1018 662
rect 1126 658 1130 662
rect 1150 658 1154 662
rect 1190 658 1194 662
rect 1214 658 1218 662
rect 1278 658 1282 662
rect 1302 658 1306 662
rect 1326 658 1330 662
rect 1334 658 1338 662
rect 1390 658 1394 662
rect 1414 658 1418 662
rect 1438 658 1442 662
rect 1486 658 1490 662
rect 1534 658 1538 662
rect 1606 658 1610 662
rect 1630 658 1634 662
rect 1638 658 1642 662
rect 1678 658 1682 662
rect 1686 658 1690 662
rect 1702 658 1706 662
rect 1750 658 1754 662
rect 1790 658 1794 662
rect 1830 658 1834 662
rect 1854 658 1858 662
rect 1870 658 1874 662
rect 1926 658 1930 662
rect 2046 658 2050 662
rect 2070 658 2074 662
rect 2094 658 2098 662
rect 2134 658 2138 662
rect 2150 658 2154 662
rect 2174 658 2178 662
rect 2222 658 2226 662
rect 2254 659 2258 663
rect 2286 658 2290 662
rect 2326 658 2330 662
rect 2366 658 2370 662
rect 2382 658 2386 662
rect 2390 658 2394 662
rect 2406 658 2410 662
rect 2446 658 2450 662
rect 2470 658 2474 662
rect 2558 659 2562 663
rect 2646 658 2650 662
rect 2678 658 2682 662
rect 2686 658 2690 662
rect 2742 659 2746 663
rect 2822 658 2826 662
rect 2886 658 2890 662
rect 2902 658 2906 662
rect 2950 658 2954 662
rect 2974 658 2978 662
rect 2990 658 2994 662
rect 3022 658 3026 662
rect 3046 658 3050 662
rect 3078 658 3082 662
rect 3118 658 3122 662
rect 3134 658 3138 662
rect 3158 658 3162 662
rect 3190 658 3194 662
rect 3214 658 3218 662
rect 3254 659 3258 663
rect 3286 658 3290 662
rect 3342 658 3346 662
rect 3358 658 3362 662
rect 3374 658 3378 662
rect 3406 658 3410 662
rect 3454 659 3458 663
rect 3526 658 3530 662
rect 54 648 58 652
rect 110 648 114 652
rect 166 648 170 652
rect 230 648 234 652
rect 270 648 274 652
rect 382 648 386 652
rect 390 648 394 652
rect 430 648 434 652
rect 454 648 458 652
rect 462 648 466 652
rect 478 648 482 652
rect 534 648 538 652
rect 582 648 586 652
rect 590 648 594 652
rect 622 648 626 652
rect 654 648 658 652
rect 734 648 738 652
rect 782 648 786 652
rect 870 648 874 652
rect 926 648 930 652
rect 958 648 962 652
rect 1030 648 1034 652
rect 1054 648 1058 652
rect 1110 648 1114 652
rect 1174 648 1178 652
rect 1230 648 1234 652
rect 1238 648 1242 652
rect 1286 648 1290 652
rect 1366 648 1370 652
rect 1398 648 1402 652
rect 1454 648 1458 652
rect 1510 648 1514 652
rect 1654 648 1658 652
rect 1694 648 1698 652
rect 1734 648 1738 652
rect 1934 648 1938 652
rect 2014 648 2018 652
rect 2054 648 2058 652
rect 2070 648 2074 652
rect 2142 648 2146 652
rect 2198 648 2202 652
rect 2398 648 2402 652
rect 2438 648 2442 652
rect 2470 648 2474 652
rect 2710 648 2714 652
rect 2838 648 2842 652
rect 2918 648 2922 652
rect 2958 648 2962 652
rect 3054 648 3058 652
rect 3134 648 3138 652
rect 3222 648 3226 652
rect 286 638 290 642
rect 710 638 714 642
rect 1214 638 1218 642
rect 1350 638 1354 642
rect 1926 638 1930 642
rect 2126 638 2130 642
rect 2462 638 2466 642
rect 2622 638 2626 642
rect 3038 638 3042 642
rect 3102 638 3106 642
rect 3206 638 3210 642
rect 3558 638 3562 642
rect 1102 628 1106 632
rect 2846 628 2850 632
rect 2926 628 2930 632
rect 606 618 610 622
rect 694 618 698 622
rect 750 618 754 622
rect 806 618 810 622
rect 1062 618 1066 622
rect 1150 618 1154 622
rect 1382 618 1386 622
rect 1414 618 1418 622
rect 1630 618 1634 622
rect 1894 618 1898 622
rect 1990 618 1994 622
rect 2134 618 2138 622
rect 2366 618 2370 622
rect 2870 618 2874 622
rect 2902 618 2906 622
rect 3046 618 3050 622
rect 3390 618 3394 622
rect 482 603 486 607
rect 489 603 493 607
rect 1514 603 1518 607
rect 1521 603 1525 607
rect 2538 603 2542 607
rect 2545 603 2549 607
rect 22 588 26 592
rect 86 588 90 592
rect 150 588 154 592
rect 182 588 186 592
rect 198 588 202 592
rect 230 588 234 592
rect 254 588 258 592
rect 398 588 402 592
rect 414 588 418 592
rect 430 588 434 592
rect 558 588 562 592
rect 622 588 626 592
rect 678 588 682 592
rect 710 588 714 592
rect 814 588 818 592
rect 878 588 882 592
rect 910 588 914 592
rect 950 588 954 592
rect 1022 588 1026 592
rect 1046 588 1050 592
rect 1166 588 1170 592
rect 1206 588 1210 592
rect 1342 588 1346 592
rect 1374 588 1378 592
rect 1478 588 1482 592
rect 1534 588 1538 592
rect 1574 588 1578 592
rect 1614 588 1618 592
rect 1638 588 1642 592
rect 1710 588 1714 592
rect 1878 588 1882 592
rect 2374 588 2378 592
rect 2566 588 2570 592
rect 2622 588 2626 592
rect 2798 588 2802 592
rect 2878 588 2882 592
rect 2990 588 2994 592
rect 3110 588 3114 592
rect 3278 588 3282 592
rect 3366 588 3370 592
rect 366 578 370 582
rect 334 568 338 572
rect 734 568 738 572
rect 1334 568 1338 572
rect 1646 568 1650 572
rect 1886 568 1890 572
rect 2366 568 2370 572
rect 2654 568 2658 572
rect 2742 568 2746 572
rect 2926 568 2930 572
rect 3094 568 3098 572
rect 3118 568 3122 572
rect 3134 568 3138 572
rect 3486 568 3490 572
rect 3534 568 3538 572
rect 270 558 274 562
rect 350 558 354 562
rect 382 558 386 562
rect 438 558 442 562
rect 494 558 498 562
rect 534 558 538 562
rect 6 548 10 552
rect 38 548 42 552
rect 70 548 74 552
rect 102 548 106 552
rect 134 548 138 552
rect 166 548 170 552
rect 214 548 218 552
rect 286 548 290 552
rect 318 548 322 552
rect 334 548 338 552
rect 366 548 370 552
rect 454 548 458 552
rect 470 548 474 552
rect 590 558 594 562
rect 718 558 722 562
rect 766 558 770 562
rect 566 548 570 552
rect 606 548 610 552
rect 654 548 658 552
rect 662 548 666 552
rect 686 548 690 552
rect 734 548 738 552
rect 782 548 786 552
rect 790 548 794 552
rect 838 558 842 562
rect 894 558 898 562
rect 918 558 922 562
rect 1030 558 1034 562
rect 1062 558 1066 562
rect 1070 558 1074 562
rect 1086 558 1090 562
rect 1118 558 1122 562
rect 854 548 858 552
rect 878 548 882 552
rect 926 548 930 552
rect 934 548 938 552
rect 958 548 962 552
rect 966 548 970 552
rect 990 548 994 552
rect 1046 548 1050 552
rect 1102 548 1106 552
rect 1110 548 1114 552
rect 1134 548 1138 552
rect 1142 548 1146 552
rect 1150 548 1154 552
rect 1182 548 1186 552
rect 1190 548 1194 552
rect 1206 548 1210 552
rect 1230 558 1234 562
rect 1294 558 1298 562
rect 1342 558 1346 562
rect 1630 558 1634 562
rect 1750 558 1754 562
rect 1782 558 1786 562
rect 1806 558 1810 562
rect 1870 558 1874 562
rect 1926 558 1930 562
rect 1950 558 1954 562
rect 1982 558 1986 562
rect 1990 558 1994 562
rect 2006 558 2010 562
rect 2046 558 2050 562
rect 2078 558 2082 562
rect 2110 558 2114 562
rect 2126 558 2130 562
rect 2142 558 2146 562
rect 2270 558 2274 562
rect 2310 558 2314 562
rect 2350 558 2354 562
rect 2606 558 2610 562
rect 2638 558 2642 562
rect 2726 558 2730 562
rect 2862 558 2866 562
rect 1246 548 1250 552
rect 1286 548 1290 552
rect 1310 548 1314 552
rect 1318 548 1322 552
rect 1342 548 1346 552
rect 1358 548 1362 552
rect 1366 548 1370 552
rect 1390 548 1394 552
rect 1406 548 1410 552
rect 1414 548 1418 552
rect 1438 548 1442 552
rect 1454 548 1458 552
rect 1462 548 1466 552
rect 1486 548 1490 552
rect 1518 548 1522 552
rect 1526 548 1530 552
rect 1550 548 1554 552
rect 1590 548 1594 552
rect 1598 548 1602 552
rect 1638 548 1642 552
rect 1662 548 1666 552
rect 1694 548 1698 552
rect 1726 548 1730 552
rect 1742 548 1746 552
rect 1758 548 1762 552
rect 1774 548 1778 552
rect 1798 548 1802 552
rect 1822 548 1826 552
rect 1878 548 1882 552
rect 1910 548 1914 552
rect 1918 548 1922 552
rect 2006 548 2010 552
rect 2014 548 2018 552
rect 2126 548 2130 552
rect 2142 548 2146 552
rect 2158 548 2162 552
rect 62 538 66 542
rect 126 538 130 542
rect 246 538 250 542
rect 286 538 290 542
rect 2198 547 2202 551
rect 2286 548 2290 552
rect 2318 548 2322 552
rect 2326 548 2330 552
rect 2358 548 2362 552
rect 2390 548 2394 552
rect 2446 548 2450 552
rect 2518 548 2522 552
rect 2582 548 2586 552
rect 2606 548 2610 552
rect 2622 548 2626 552
rect 2646 548 2650 552
rect 2670 548 2674 552
rect 2686 548 2690 552
rect 2702 548 2706 552
rect 2710 548 2714 552
rect 2734 548 2738 552
rect 2758 548 2762 552
rect 2798 548 2802 552
rect 2854 548 2858 552
rect 2878 548 2882 552
rect 2974 558 2978 562
rect 3006 558 3010 562
rect 3014 558 3018 562
rect 3054 558 3058 562
rect 3102 558 3106 562
rect 3246 558 3250 562
rect 3390 558 3394 562
rect 2918 548 2922 552
rect 2926 548 2930 552
rect 2958 548 2962 552
rect 2966 548 2970 552
rect 2990 548 2994 552
rect 3006 548 3010 552
rect 3030 548 3034 552
rect 3070 548 3074 552
rect 3118 548 3122 552
rect 3166 548 3170 552
rect 3190 548 3194 552
rect 3230 548 3234 552
rect 3286 548 3290 552
rect 3326 548 3330 552
rect 3342 548 3346 552
rect 3422 547 3426 551
rect 3494 548 3498 552
rect 3518 548 3522 552
rect 326 538 330 542
rect 358 538 362 542
rect 422 538 426 542
rect 438 538 442 542
rect 478 538 482 542
rect 518 538 522 542
rect 566 538 570 542
rect 614 538 618 542
rect 638 538 642 542
rect 742 538 746 542
rect 750 538 754 542
rect 798 538 802 542
rect 806 538 810 542
rect 870 538 874 542
rect 902 538 906 542
rect 1014 538 1018 542
rect 1030 538 1034 542
rect 1094 538 1098 542
rect 1198 538 1202 542
rect 1686 538 1690 542
rect 1718 538 1722 542
rect 1798 538 1802 542
rect 1830 538 1834 542
rect 1846 538 1850 542
rect 1902 538 1906 542
rect 1934 538 1938 542
rect 1958 538 1962 542
rect 2014 538 2018 542
rect 2062 538 2066 542
rect 2134 538 2138 542
rect 2166 538 2170 542
rect 2214 538 2218 542
rect 2294 538 2298 542
rect 2310 538 2314 542
rect 2478 538 2482 542
rect 2494 538 2498 542
rect 2510 538 2514 542
rect 2550 538 2554 542
rect 2590 538 2594 542
rect 2630 538 2634 542
rect 2678 538 2682 542
rect 2694 538 2698 542
rect 2750 538 2754 542
rect 2814 538 2818 542
rect 2838 538 2842 542
rect 2870 538 2874 542
rect 2950 538 2954 542
rect 2982 538 2986 542
rect 3030 538 3034 542
rect 3078 538 3082 542
rect 3150 538 3154 542
rect 3182 538 3186 542
rect 3190 538 3194 542
rect 3222 538 3226 542
rect 3286 538 3290 542
rect 3302 538 3306 542
rect 3374 538 3378 542
rect 3438 538 3442 542
rect 3454 538 3458 542
rect 3510 538 3514 542
rect 3542 538 3546 542
rect 206 528 210 532
rect 390 528 394 532
rect 406 528 410 532
rect 646 528 650 532
rect 702 528 706 532
rect 990 528 994 532
rect 1270 528 1274 532
rect 1710 528 1714 532
rect 1862 528 1866 532
rect 2054 528 2058 532
rect 2086 528 2090 532
rect 2102 528 2106 532
rect 2270 528 2274 532
rect 2390 528 2394 532
rect 2494 528 2498 532
rect 2526 528 2530 532
rect 2574 528 2578 532
rect 2710 528 2714 532
rect 2782 528 2786 532
rect 2806 528 2810 532
rect 2902 528 2906 532
rect 2942 528 2946 532
rect 3094 528 3098 532
rect 3166 528 3170 532
rect 3182 528 3186 532
rect 3214 528 3218 532
rect 3326 528 3330 532
rect 3342 528 3346 532
rect 22 518 26 522
rect 230 518 234 522
rect 270 518 274 522
rect 1430 518 1434 522
rect 1614 518 1618 522
rect 1854 518 1858 522
rect 1950 518 1954 522
rect 1982 518 1986 522
rect 2342 518 2346 522
rect 2662 518 2666 522
rect 2774 518 2778 522
rect 3206 518 3210 522
rect 3246 518 3250 522
rect 3382 518 3386 522
rect 3558 518 3562 522
rect 994 503 998 507
rect 1001 503 1005 507
rect 2026 503 2030 507
rect 2033 503 2037 507
rect 3042 503 3046 507
rect 3049 503 3053 507
rect 30 488 34 492
rect 62 488 66 492
rect 78 488 82 492
rect 110 488 114 492
rect 142 488 146 492
rect 222 488 226 492
rect 254 488 258 492
rect 318 488 322 492
rect 342 488 346 492
rect 414 488 418 492
rect 478 488 482 492
rect 598 488 602 492
rect 638 488 642 492
rect 654 488 658 492
rect 694 488 698 492
rect 806 488 810 492
rect 822 488 826 492
rect 846 488 850 492
rect 862 488 866 492
rect 934 488 938 492
rect 982 488 986 492
rect 1046 488 1050 492
rect 1094 488 1098 492
rect 1222 488 1226 492
rect 1270 488 1274 492
rect 1318 488 1322 492
rect 1438 488 1442 492
rect 1582 488 1586 492
rect 1758 488 1762 492
rect 1838 488 1842 492
rect 2006 488 2010 492
rect 2102 488 2106 492
rect 2262 488 2266 492
rect 2310 488 2314 492
rect 2374 488 2378 492
rect 2406 488 2410 492
rect 2430 488 2434 492
rect 2486 488 2490 492
rect 2518 488 2522 492
rect 2526 488 2530 492
rect 2606 488 2610 492
rect 2630 488 2634 492
rect 2702 488 2706 492
rect 2742 488 2746 492
rect 2782 488 2786 492
rect 2830 488 2834 492
rect 2910 488 2914 492
rect 2934 488 2938 492
rect 2998 488 3002 492
rect 3118 488 3122 492
rect 3190 488 3194 492
rect 3198 488 3202 492
rect 3350 488 3354 492
rect 3534 488 3538 492
rect 3550 488 3554 492
rect 86 478 90 482
rect 262 478 266 482
rect 310 478 314 482
rect 646 478 650 482
rect 710 478 714 482
rect 750 478 754 482
rect 854 478 858 482
rect 926 478 930 482
rect 942 478 946 482
rect 990 478 994 482
rect 1430 478 1434 482
rect 1550 478 1554 482
rect 1566 478 1570 482
rect 1670 478 1674 482
rect 1678 478 1682 482
rect 1878 478 1882 482
rect 38 468 42 472
rect 150 468 154 472
rect 174 468 178 472
rect 206 468 210 472
rect 222 468 226 472
rect 302 468 306 472
rect 326 468 330 472
rect 350 468 354 472
rect 366 468 370 472
rect 398 468 402 472
rect 406 468 410 472
rect 510 468 514 472
rect 558 468 562 472
rect 598 468 602 472
rect 614 468 618 472
rect 622 468 626 472
rect 662 468 666 472
rect 686 468 690 472
rect 758 468 762 472
rect 782 468 786 472
rect 830 468 834 472
rect 886 468 890 472
rect 46 458 50 462
rect 94 458 98 462
rect 126 458 130 462
rect 166 458 170 462
rect 206 458 210 462
rect 230 458 234 462
rect 278 458 282 462
rect 390 458 394 462
rect 430 458 434 462
rect 462 458 466 462
rect 534 458 538 462
rect 550 458 554 462
rect 558 458 562 462
rect 582 458 586 462
rect 726 458 730 462
rect 782 458 786 462
rect 838 458 842 462
rect 878 458 882 462
rect 910 468 914 472
rect 1038 468 1042 472
rect 1062 468 1066 472
rect 1070 468 1074 472
rect 1142 468 1146 472
rect 1190 468 1194 472
rect 1342 468 1346 472
rect 1390 468 1394 472
rect 1398 468 1402 472
rect 1446 468 1450 472
rect 1486 468 1490 472
rect 1518 468 1522 472
rect 1574 468 1578 472
rect 1606 468 1610 472
rect 1614 468 1618 472
rect 1630 468 1634 472
rect 1654 468 1658 472
rect 1694 468 1698 472
rect 1710 468 1714 472
rect 1798 468 1802 472
rect 1846 468 1850 472
rect 2054 478 2058 482
rect 2110 478 2114 482
rect 2238 478 2242 482
rect 2558 478 2562 482
rect 2638 478 2642 482
rect 2654 478 2658 482
rect 2662 478 2666 482
rect 2670 478 2674 482
rect 2726 478 2730 482
rect 2734 478 2738 482
rect 2774 478 2778 482
rect 2838 478 2842 482
rect 2862 478 2866 482
rect 2878 478 2882 482
rect 3022 478 3026 482
rect 3110 478 3114 482
rect 3222 478 3226 482
rect 3254 478 3258 482
rect 3342 478 3346 482
rect 3414 478 3418 482
rect 1894 468 1898 472
rect 1934 468 1938 472
rect 1982 468 1986 472
rect 1998 468 2002 472
rect 2014 468 2018 472
rect 2054 468 2058 472
rect 2086 468 2090 472
rect 2142 468 2146 472
rect 2174 468 2178 472
rect 2190 468 2194 472
rect 2230 468 2234 472
rect 2254 468 2258 472
rect 2302 468 2306 472
rect 2334 468 2338 472
rect 2342 468 2346 472
rect 2398 468 2402 472
rect 2422 468 2426 472
rect 2454 468 2458 472
rect 2494 468 2498 472
rect 2582 468 2586 472
rect 2598 468 2602 472
rect 2622 468 2626 472
rect 2766 468 2770 472
rect 2790 468 2794 472
rect 2806 468 2810 472
rect 2886 468 2890 472
rect 2926 468 2930 472
rect 2958 468 2962 472
rect 2974 468 2978 472
rect 2990 468 2994 472
rect 3038 468 3042 472
rect 3070 468 3074 472
rect 3094 468 3098 472
rect 3150 468 3154 472
rect 3158 468 3162 472
rect 3166 468 3170 472
rect 3238 468 3242 472
rect 3270 468 3274 472
rect 3294 468 3298 472
rect 3310 468 3314 472
rect 3326 468 3330 472
rect 3374 468 3378 472
rect 3430 468 3434 472
rect 3454 468 3458 472
rect 3542 468 3546 472
rect 902 458 906 462
rect 958 458 962 462
rect 974 458 978 462
rect 990 458 994 462
rect 1030 458 1034 462
rect 1070 458 1074 462
rect 1102 458 1106 462
rect 1110 458 1114 462
rect 1134 458 1138 462
rect 1150 458 1154 462
rect 1158 458 1162 462
rect 1182 458 1186 462
rect 1198 458 1202 462
rect 1206 458 1210 462
rect 1230 458 1234 462
rect 1246 458 1250 462
rect 1254 458 1258 462
rect 1278 458 1282 462
rect 1294 458 1298 462
rect 1302 458 1306 462
rect 1326 458 1330 462
rect 1406 458 1410 462
rect 1430 458 1434 462
rect 1446 458 1450 462
rect 1478 458 1482 462
rect 1494 458 1498 462
rect 1534 458 1538 462
rect 1598 458 1602 462
rect 1622 458 1626 462
rect 1646 458 1650 462
rect 1662 458 1666 462
rect 1686 458 1690 462
rect 1710 458 1714 462
rect 1718 458 1722 462
rect 1782 458 1786 462
rect 1806 458 1810 462
rect 1854 458 1858 462
rect 1862 458 1866 462
rect 1918 458 1922 462
rect 1974 458 1978 462
rect 1990 458 1994 462
rect 2022 458 2026 462
rect 2062 458 2066 462
rect 2078 458 2082 462
rect 2142 458 2146 462
rect 2174 458 2178 462
rect 2182 458 2186 462
rect 2246 458 2250 462
rect 2302 458 2306 462
rect 2326 458 2330 462
rect 2350 458 2354 462
rect 2374 458 2378 462
rect 2390 458 2394 462
rect 2446 458 2450 462
rect 2502 458 2506 462
rect 2598 458 2602 462
rect 2614 458 2618 462
rect 2646 458 2650 462
rect 2686 458 2690 462
rect 2702 458 2706 462
rect 2758 458 2762 462
rect 2798 458 2802 462
rect 2854 458 2858 462
rect 2878 458 2882 462
rect 2950 458 2954 462
rect 2982 458 2986 462
rect 3054 458 3058 462
rect 3086 458 3090 462
rect 3118 458 3122 462
rect 3142 458 3146 462
rect 3174 458 3178 462
rect 3246 458 3250 462
rect 3262 458 3266 462
rect 3278 458 3282 462
rect 3302 458 3306 462
rect 3318 458 3322 462
rect 3366 458 3370 462
rect 3398 458 3402 462
rect 3438 458 3442 462
rect 3470 459 3474 463
rect 182 448 186 452
rect 222 448 226 452
rect 254 448 258 452
rect 262 448 266 452
rect 342 448 346 452
rect 366 448 370 452
rect 422 448 426 452
rect 526 448 530 452
rect 534 448 538 452
rect 566 448 570 452
rect 598 448 602 452
rect 638 448 642 452
rect 678 448 682 452
rect 686 448 690 452
rect 702 448 706 452
rect 750 448 754 452
rect 758 448 762 452
rect 774 448 778 452
rect 806 448 810 452
rect 814 448 818 452
rect 862 448 866 452
rect 918 448 922 452
rect 942 448 946 452
rect 1014 448 1018 452
rect 1046 448 1050 452
rect 1094 448 1098 452
rect 1422 448 1426 452
rect 1510 448 1514 452
rect 1582 448 1586 452
rect 1638 448 1642 452
rect 1734 448 1738 452
rect 1758 448 1762 452
rect 1790 448 1794 452
rect 1822 448 1826 452
rect 1926 448 1930 452
rect 1950 448 1954 452
rect 1958 448 1962 452
rect 1974 448 1978 452
rect 2054 448 2058 452
rect 2118 448 2122 452
rect 2134 448 2138 452
rect 2150 448 2154 452
rect 2278 448 2282 452
rect 2310 448 2314 452
rect 2366 448 2370 452
rect 2374 448 2378 452
rect 2406 448 2410 452
rect 2430 448 2434 452
rect 2486 448 2490 452
rect 2518 448 2522 452
rect 2526 448 2530 452
rect 2694 448 2698 452
rect 2742 448 2746 452
rect 2830 448 2834 452
rect 2902 448 2906 452
rect 2910 448 2914 452
rect 2934 448 2938 452
rect 2966 448 2970 452
rect 2998 448 3002 452
rect 3118 448 3122 452
rect 3190 448 3194 452
rect 3198 448 3202 452
rect 3286 448 3290 452
rect 3382 448 3386 452
rect 3398 448 3402 452
rect 1774 438 1778 442
rect 1910 438 1914 442
rect 2166 438 2170 442
rect 2710 438 2714 442
rect 518 428 522 432
rect 3078 428 3082 432
rect 30 418 34 422
rect 446 418 450 422
rect 1374 418 1378 422
rect 1462 418 1466 422
rect 1766 418 1770 422
rect 1918 418 1922 422
rect 1942 418 1946 422
rect 2206 418 2210 422
rect 2678 418 2682 422
rect 2846 418 2850 422
rect 482 403 486 407
rect 489 403 493 407
rect 1514 403 1518 407
rect 1521 403 1525 407
rect 2538 403 2542 407
rect 2545 403 2549 407
rect 22 388 26 392
rect 54 388 58 392
rect 86 388 90 392
rect 118 388 122 392
rect 150 388 154 392
rect 206 388 210 392
rect 278 388 282 392
rect 334 388 338 392
rect 366 388 370 392
rect 382 388 386 392
rect 414 388 418 392
rect 470 388 474 392
rect 526 388 530 392
rect 606 388 610 392
rect 678 388 682 392
rect 694 388 698 392
rect 790 388 794 392
rect 838 388 842 392
rect 934 388 938 392
rect 966 388 970 392
rect 982 388 986 392
rect 1086 388 1090 392
rect 1126 388 1130 392
rect 1174 388 1178 392
rect 1230 388 1234 392
rect 1302 388 1306 392
rect 1342 388 1346 392
rect 1430 388 1434 392
rect 1478 388 1482 392
rect 1638 388 1642 392
rect 1734 388 1738 392
rect 1774 388 1778 392
rect 1822 388 1826 392
rect 2014 388 2018 392
rect 2134 388 2138 392
rect 2230 388 2234 392
rect 2302 388 2306 392
rect 2350 388 2354 392
rect 2454 388 2458 392
rect 2494 388 2498 392
rect 2574 388 2578 392
rect 2590 388 2594 392
rect 2654 388 2658 392
rect 2710 388 2714 392
rect 2750 388 2754 392
rect 2790 388 2794 392
rect 2902 388 2906 392
rect 3030 388 3034 392
rect 3142 388 3146 392
rect 3174 388 3178 392
rect 3278 388 3282 392
rect 3366 388 3370 392
rect 3502 388 3506 392
rect 2478 378 2482 382
rect 3486 378 3490 382
rect 558 368 562 372
rect 1678 368 1682 372
rect 2142 368 2146 372
rect 2710 368 2714 372
rect 2718 368 2722 372
rect 2854 368 2858 372
rect 3022 368 3026 372
rect 3102 368 3106 372
rect 3406 368 3410 372
rect 222 358 226 362
rect 310 358 314 362
rect 6 348 10 352
rect 38 348 42 352
rect 70 348 74 352
rect 102 348 106 352
rect 134 348 138 352
rect 158 348 162 352
rect 166 348 170 352
rect 206 348 210 352
rect 230 348 234 352
rect 262 348 266 352
rect 350 358 354 362
rect 398 358 402 362
rect 494 358 498 362
rect 542 358 546 362
rect 334 348 338 352
rect 366 348 370 352
rect 414 348 418 352
rect 454 348 458 352
rect 478 348 482 352
rect 502 348 506 352
rect 526 348 530 352
rect 566 358 570 362
rect 582 348 586 352
rect 606 348 610 352
rect 630 358 634 362
rect 662 358 666 362
rect 758 358 762 362
rect 862 358 866 362
rect 870 358 874 362
rect 886 358 890 362
rect 918 358 922 362
rect 950 358 954 362
rect 1038 358 1042 362
rect 1254 358 1258 362
rect 646 348 650 352
rect 678 348 682 352
rect 694 348 698 352
rect 742 348 746 352
rect 758 348 762 352
rect 766 348 770 352
rect 774 348 778 352
rect 798 348 802 352
rect 814 348 818 352
rect 822 348 826 352
rect 846 348 850 352
rect 918 348 922 352
rect 934 348 938 352
rect 966 348 970 352
rect 1006 348 1010 352
rect 1022 348 1026 352
rect 1046 348 1050 352
rect 1054 348 1058 352
rect 1070 348 1074 352
rect 1094 348 1098 352
rect 1110 348 1114 352
rect 1118 348 1122 352
rect 1142 348 1146 352
rect 1158 348 1162 352
rect 1166 348 1170 352
rect 1190 348 1194 352
rect 1198 348 1202 352
rect 1214 348 1218 352
rect 1238 348 1242 352
rect 1278 348 1282 352
rect 1286 348 1290 352
rect 1310 348 1314 352
rect 1326 348 1330 352
rect 1334 348 1338 352
rect 1358 348 1362 352
rect 1366 348 1370 352
rect 1398 348 1402 352
rect 1486 348 1490 352
rect 1606 348 1610 352
rect 1622 348 1626 352
rect 1662 358 1666 362
rect 1894 358 1898 362
rect 1942 358 1946 362
rect 1974 358 1978 362
rect 2006 358 2010 362
rect 2046 358 2050 362
rect 2078 358 2082 362
rect 2158 358 2162 362
rect 2214 358 2218 362
rect 2246 358 2250 362
rect 2334 358 2338 362
rect 2358 358 2362 362
rect 2414 358 2418 362
rect 2526 358 2530 362
rect 2606 358 2610 362
rect 2702 358 2706 362
rect 2734 358 2738 362
rect 2806 358 2810 362
rect 2814 358 2818 362
rect 2870 358 2874 362
rect 2958 358 2962 362
rect 3046 358 3050 362
rect 3158 358 3162 362
rect 3190 358 3194 362
rect 3222 358 3226 362
rect 3246 358 3250 362
rect 3270 358 3274 362
rect 3318 358 3322 362
rect 1678 348 1682 352
rect 1718 348 1722 352
rect 1742 348 1746 352
rect 1750 348 1754 352
rect 1782 348 1786 352
rect 1814 348 1818 352
rect 1846 348 1850 352
rect 1854 348 1858 352
rect 1902 348 1906 352
rect 1982 348 1986 352
rect 2006 348 2010 352
rect 2030 348 2034 352
rect 2062 348 2066 352
rect 2102 348 2106 352
rect 2150 348 2154 352
rect 2174 348 2178 352
rect 2182 348 2186 352
rect 2190 348 2194 352
rect 2206 348 2210 352
rect 2246 348 2250 352
rect 2278 348 2282 352
rect 2318 348 2322 352
rect 2366 348 2370 352
rect 2374 348 2378 352
rect 2382 348 2386 352
rect 2406 348 2410 352
rect 2422 348 2426 352
rect 2510 348 2514 352
rect 2518 348 2522 352
rect 2550 348 2554 352
rect 2590 348 2594 352
rect 2638 348 2642 352
rect 182 338 186 342
rect 198 338 202 342
rect 246 338 250 342
rect 286 338 290 342
rect 342 338 346 342
rect 374 338 378 342
rect 534 338 538 342
rect 542 338 546 342
rect 590 338 594 342
rect 598 338 602 342
rect 654 338 658 342
rect 686 338 690 342
rect 878 338 882 342
rect 894 338 898 342
rect 910 338 914 342
rect 942 338 946 342
rect 974 338 978 342
rect 1270 338 1274 342
rect 1398 338 1402 342
rect 1406 338 1410 342
rect 1446 338 1450 342
rect 1470 338 1474 342
rect 1526 338 1530 342
rect 1542 338 1546 342
rect 1550 338 1554 342
rect 1598 338 1602 342
rect 1630 338 1634 342
rect 1686 338 1690 342
rect 1710 338 1714 342
rect 1750 338 1754 342
rect 1790 338 1794 342
rect 1822 338 1826 342
rect 1838 338 1842 342
rect 1878 338 1882 342
rect 1926 338 1930 342
rect 1950 338 1954 342
rect 1966 338 1970 342
rect 2022 338 2026 342
rect 2070 338 2074 342
rect 2078 338 2082 342
rect 2094 338 2098 342
rect 2110 338 2114 342
rect 2190 338 2194 342
rect 2222 338 2226 342
rect 2310 338 2314 342
rect 2326 338 2330 342
rect 2382 338 2386 342
rect 2390 338 2394 342
rect 2430 338 2434 342
rect 2462 338 2466 342
rect 2470 338 2474 342
rect 2502 338 2506 342
rect 2558 338 2562 342
rect 2582 338 2586 342
rect 2630 338 2634 342
rect 2678 348 2682 352
rect 2710 348 2714 352
rect 2750 348 2754 352
rect 2814 348 2818 352
rect 2830 348 2834 352
rect 2854 348 2858 352
rect 2878 348 2882 352
rect 2942 348 2946 352
rect 3006 348 3010 352
rect 3030 348 3034 352
rect 3062 348 3066 352
rect 3078 348 3082 352
rect 3094 348 3098 352
rect 3126 348 3130 352
rect 3142 348 3146 352
rect 3166 348 3170 352
rect 3206 348 3210 352
rect 3286 348 3290 352
rect 3350 348 3354 352
rect 3374 348 3378 352
rect 3382 348 3386 352
rect 3414 348 3418 352
rect 3430 348 3434 352
rect 3446 348 3450 352
rect 2654 338 2658 342
rect 2670 338 2674 342
rect 2782 338 2786 342
rect 2838 338 2842 342
rect 2846 338 2850 342
rect 2886 338 2890 342
rect 2910 338 2914 342
rect 2934 338 2938 342
rect 2998 338 3002 342
rect 3046 338 3050 342
rect 3070 338 3074 342
rect 3086 338 3090 342
rect 3118 338 3122 342
rect 3134 338 3138 342
rect 3166 338 3170 342
rect 3198 338 3202 342
rect 3214 338 3218 342
rect 3230 338 3234 342
rect 3246 338 3250 342
rect 3262 338 3266 342
rect 3286 338 3290 342
rect 3318 338 3322 342
rect 3334 338 3338 342
rect 3382 338 3386 342
rect 3406 338 3410 342
rect 3438 338 3442 342
rect 3470 348 3474 352
rect 3510 348 3514 352
rect 3518 348 3522 352
rect 3534 348 3538 352
rect 390 328 394 332
rect 438 328 442 332
rect 710 328 714 332
rect 726 328 730 332
rect 990 328 994 332
rect 1374 328 1378 332
rect 1462 328 1466 332
rect 1606 328 1610 332
rect 1694 328 1698 332
rect 1726 328 1730 332
rect 1774 328 1778 332
rect 1806 328 1810 332
rect 1870 328 1874 332
rect 1918 328 1922 332
rect 1998 328 2002 332
rect 2126 328 2130 332
rect 2166 328 2170 332
rect 2270 328 2274 332
rect 2302 328 2306 332
rect 2342 328 2346 332
rect 2438 328 2442 332
rect 2446 328 2450 332
rect 2486 328 2490 332
rect 2574 328 2578 332
rect 2614 328 2618 332
rect 2622 328 2626 332
rect 2686 328 2690 332
rect 2774 328 2778 332
rect 2902 328 2906 332
rect 2910 328 2914 332
rect 2966 328 2970 332
rect 3102 328 3106 332
rect 3310 328 3314 332
rect 3350 328 3354 332
rect 3358 328 3362 332
rect 3422 328 3426 332
rect 3470 328 3474 332
rect 3494 328 3498 332
rect 3542 328 3546 332
rect 718 318 722 322
rect 1262 318 1266 322
rect 1414 318 1418 322
rect 1454 318 1458 322
rect 1518 318 1522 322
rect 1582 318 1586 322
rect 1702 318 1706 322
rect 1798 318 1802 322
rect 1862 318 1866 322
rect 1894 318 1898 322
rect 1910 318 1914 322
rect 1942 318 1946 322
rect 2006 318 2010 322
rect 2118 318 2122 322
rect 2958 318 2962 322
rect 2990 318 2994 322
rect 3254 318 3258 322
rect 3302 318 3306 322
rect 994 303 998 307
rect 1001 303 1005 307
rect 2026 303 2030 307
rect 2033 303 2037 307
rect 3042 303 3046 307
rect 3049 303 3053 307
rect 22 288 26 292
rect 174 288 178 292
rect 206 288 210 292
rect 230 288 234 292
rect 254 288 258 292
rect 350 288 354 292
rect 358 288 362 292
rect 382 288 386 292
rect 398 288 402 292
rect 446 288 450 292
rect 494 288 498 292
rect 534 288 538 292
rect 542 288 546 292
rect 574 288 578 292
rect 622 288 626 292
rect 694 288 698 292
rect 758 288 762 292
rect 782 288 786 292
rect 838 288 842 292
rect 870 288 874 292
rect 950 288 954 292
rect 1030 288 1034 292
rect 1062 288 1066 292
rect 1222 288 1226 292
rect 1246 288 1250 292
rect 1350 288 1354 292
rect 1366 288 1370 292
rect 1390 288 1394 292
rect 1422 288 1426 292
rect 1694 288 1698 292
rect 1750 288 1754 292
rect 1790 288 1794 292
rect 1814 288 1818 292
rect 1830 288 1834 292
rect 1942 288 1946 292
rect 2254 288 2258 292
rect 2334 288 2338 292
rect 2390 288 2394 292
rect 2470 288 2474 292
rect 2486 288 2490 292
rect 2526 288 2530 292
rect 2590 288 2594 292
rect 2750 288 2754 292
rect 2806 288 2810 292
rect 2870 288 2874 292
rect 2894 288 2898 292
rect 2974 288 2978 292
rect 3014 288 3018 292
rect 3070 288 3074 292
rect 3094 288 3098 292
rect 3222 288 3226 292
rect 3358 288 3362 292
rect 3510 288 3514 292
rect 86 278 90 282
rect 390 278 394 282
rect 582 278 586 282
rect 854 278 858 282
rect 1022 278 1026 282
rect 1142 278 1146 282
rect 1374 278 1378 282
rect 1382 278 1386 282
rect 1430 278 1434 282
rect 1438 278 1442 282
rect 1454 278 1458 282
rect 1494 278 1498 282
rect 1526 278 1530 282
rect 1606 278 1610 282
rect 1710 278 1714 282
rect 1758 278 1762 282
rect 1822 278 1826 282
rect 1862 278 1866 282
rect 1966 278 1970 282
rect 2014 278 2018 282
rect 2086 278 2090 282
rect 2286 278 2290 282
rect 2326 278 2330 282
rect 2382 278 2386 282
rect 2438 278 2442 282
rect 2518 278 2522 282
rect 2630 278 2634 282
rect 2678 278 2682 282
rect 2686 278 2690 282
rect 2702 278 2706 282
rect 2814 278 2818 282
rect 2918 278 2922 282
rect 2926 278 2930 282
rect 2966 278 2970 282
rect 3062 278 3066 282
rect 3078 278 3082 282
rect 3142 278 3146 282
rect 3182 278 3186 282
rect 62 268 66 272
rect 222 268 226 272
rect 238 268 242 272
rect 270 268 274 272
rect 318 268 322 272
rect 6 258 10 262
rect 30 258 34 262
rect 70 258 74 262
rect 134 258 138 262
rect 166 258 170 262
rect 190 258 194 262
rect 262 258 266 262
rect 278 258 282 262
rect 286 258 290 262
rect 318 258 322 262
rect 374 268 378 272
rect 414 268 418 272
rect 470 268 474 272
rect 510 268 514 272
rect 566 268 570 272
rect 590 268 594 272
rect 614 268 618 272
rect 662 268 666 272
rect 670 268 674 272
rect 686 268 690 272
rect 718 268 722 272
rect 750 268 754 272
rect 774 268 778 272
rect 806 268 810 272
rect 814 268 818 272
rect 862 268 866 272
rect 894 268 898 272
rect 910 268 914 272
rect 926 268 930 272
rect 934 268 938 272
rect 950 268 954 272
rect 1014 268 1018 272
rect 1038 268 1042 272
rect 1102 268 1106 272
rect 1110 268 1114 272
rect 1126 268 1130 272
rect 1166 268 1170 272
rect 1174 268 1178 272
rect 1270 268 1274 272
rect 1278 268 1282 272
rect 1326 268 1330 272
rect 1334 268 1338 272
rect 1414 268 1418 272
rect 1454 268 1458 272
rect 1478 268 1482 272
rect 1550 268 1554 272
rect 1574 268 1578 272
rect 1582 268 1586 272
rect 1606 268 1610 272
rect 1646 268 1650 272
rect 1678 268 1682 272
rect 1686 268 1690 272
rect 1726 268 1730 272
rect 1742 268 1746 272
rect 1766 268 1770 272
rect 1806 268 1810 272
rect 1854 268 1858 272
rect 1878 268 1882 272
rect 1902 268 1906 272
rect 1918 268 1922 272
rect 1926 268 1930 272
rect 1950 268 1954 272
rect 2078 268 2082 272
rect 2102 268 2106 272
rect 2126 268 2130 272
rect 334 258 338 262
rect 430 258 434 262
rect 454 258 458 262
rect 462 258 466 262
rect 510 258 514 262
rect 558 258 562 262
rect 630 258 634 262
rect 654 258 658 262
rect 694 258 698 262
rect 710 258 714 262
rect 726 258 730 262
rect 742 258 746 262
rect 798 258 802 262
rect 814 258 818 262
rect 894 258 898 262
rect 926 258 930 262
rect 990 258 994 262
rect 1038 258 1042 262
rect 1046 258 1050 262
rect 1094 258 1098 262
rect 1118 258 1122 262
rect 1158 258 1162 262
rect 1166 258 1170 262
rect 1206 258 1210 262
rect 1230 258 1234 262
rect 1238 258 1242 262
rect 1270 258 1274 262
rect 1318 258 1322 262
rect 1398 258 1402 262
rect 1406 258 1410 262
rect 1454 258 1458 262
rect 1470 258 1474 262
rect 1486 258 1490 262
rect 1542 258 1546 262
rect 1550 258 1554 262
rect 2150 268 2154 272
rect 2198 268 2202 272
rect 2206 268 2210 272
rect 2222 268 2226 272
rect 2270 268 2274 272
rect 2294 268 2298 272
rect 2342 268 2346 272
rect 2486 268 2490 272
rect 2502 268 2506 272
rect 2534 268 2538 272
rect 2566 268 2570 272
rect 2622 268 2626 272
rect 2638 268 2642 272
rect 2662 268 2666 272
rect 2710 268 2714 272
rect 2734 268 2738 272
rect 2782 268 2786 272
rect 2798 268 2802 272
rect 2814 268 2818 272
rect 2846 268 2850 272
rect 2854 268 2858 272
rect 2878 268 2882 272
rect 2910 268 2914 272
rect 2934 268 2938 272
rect 2950 268 2954 272
rect 2990 268 2994 272
rect 3078 268 3082 272
rect 3110 268 3114 272
rect 3126 268 3130 272
rect 3166 268 3170 272
rect 3206 268 3210 272
rect 3238 268 3242 272
rect 3254 268 3258 272
rect 3262 268 3266 272
rect 3278 278 3282 282
rect 3414 278 3418 282
rect 3326 268 3330 272
rect 3390 268 3394 272
rect 3406 268 3410 272
rect 3438 268 3442 272
rect 3454 268 3458 272
rect 3470 268 3474 272
rect 3518 268 3522 272
rect 3542 278 3546 282
rect 1638 258 1642 262
rect 1670 258 1674 262
rect 1702 258 1706 262
rect 1726 258 1730 262
rect 1734 258 1738 262
rect 1774 258 1778 262
rect 1798 258 1802 262
rect 1846 258 1850 262
rect 1870 258 1874 262
rect 1886 258 1890 262
rect 1910 258 1914 262
rect 1998 258 2002 262
rect 2030 258 2034 262
rect 2054 258 2058 262
rect 2070 258 2074 262
rect 2094 258 2098 262
rect 2110 258 2114 262
rect 2134 258 2138 262
rect 2142 258 2146 262
rect 2238 258 2242 262
rect 2262 258 2266 262
rect 2302 258 2306 262
rect 2318 258 2322 262
rect 2350 258 2354 262
rect 2358 258 2362 262
rect 2398 258 2402 262
rect 2406 258 2410 262
rect 2454 258 2458 262
rect 2478 258 2482 262
rect 2510 258 2514 262
rect 2542 258 2546 262
rect 2566 258 2570 262
rect 2614 258 2618 262
rect 2790 258 2794 262
rect 2894 258 2898 262
rect 2942 258 2946 262
rect 2982 258 2986 262
rect 2998 258 3002 262
rect 3022 258 3026 262
rect 3062 258 3066 262
rect 3126 258 3130 262
rect 3166 258 3170 262
rect 3198 258 3202 262
rect 3214 258 3218 262
rect 3294 258 3298 262
rect 3398 258 3402 262
rect 3430 258 3434 262
rect 3494 258 3498 262
rect 3558 258 3562 262
rect 110 248 114 252
rect 182 248 186 252
rect 246 248 250 252
rect 262 248 266 252
rect 294 248 298 252
rect 350 248 354 252
rect 398 248 402 252
rect 534 248 538 252
rect 542 248 546 252
rect 606 248 610 252
rect 630 248 634 252
rect 638 248 642 252
rect 694 248 698 252
rect 726 248 730 252
rect 758 248 762 252
rect 782 248 786 252
rect 838 248 842 252
rect 846 248 850 252
rect 870 248 874 252
rect 902 248 906 252
rect 966 248 970 252
rect 1078 248 1082 252
rect 1142 248 1146 252
rect 1190 248 1194 252
rect 1246 248 1250 252
rect 1294 248 1298 252
rect 1574 248 1578 252
rect 1598 248 1602 252
rect 1654 248 1658 252
rect 1670 248 1674 252
rect 1830 248 1834 252
rect 1894 248 1898 252
rect 1942 248 1946 252
rect 2006 248 2010 252
rect 2054 248 2058 252
rect 2070 248 2074 252
rect 2118 248 2122 252
rect 2206 248 2210 252
rect 2254 248 2258 252
rect 2318 248 2322 252
rect 2438 248 2442 252
rect 2470 248 2474 252
rect 2598 248 2602 252
rect 2726 248 2730 252
rect 2822 248 2826 252
rect 2870 248 2874 252
rect 2958 248 2962 252
rect 3102 248 3106 252
rect 3150 248 3154 252
rect 3222 248 3226 252
rect 3318 248 3322 252
rect 3382 248 3386 252
rect 3502 248 3506 252
rect 318 238 322 242
rect 742 238 746 242
rect 1350 238 1354 242
rect 1542 238 1546 242
rect 1974 238 1978 242
rect 1982 238 1986 242
rect 1990 238 1994 242
rect 2222 238 2226 242
rect 2286 238 2290 242
rect 3486 238 3490 242
rect 1958 228 1962 232
rect 2038 228 2042 232
rect 2718 228 2722 232
rect 598 218 602 222
rect 1318 218 1322 222
rect 1502 218 1506 222
rect 1534 218 1538 222
rect 1590 218 1594 222
rect 1638 218 1642 222
rect 2374 218 2378 222
rect 2422 218 2426 222
rect 3022 218 3026 222
rect 3302 218 3306 222
rect 3342 218 3346 222
rect 3462 218 3466 222
rect 482 203 486 207
rect 489 203 493 207
rect 1514 203 1518 207
rect 1521 203 1525 207
rect 2538 203 2542 207
rect 2545 203 2549 207
rect 110 188 114 192
rect 150 188 154 192
rect 182 188 186 192
rect 358 188 362 192
rect 510 188 514 192
rect 534 188 538 192
rect 614 188 618 192
rect 750 188 754 192
rect 790 188 794 192
rect 830 188 834 192
rect 886 188 890 192
rect 918 188 922 192
rect 966 188 970 192
rect 1030 188 1034 192
rect 1070 188 1074 192
rect 1126 188 1130 192
rect 1174 188 1178 192
rect 1318 188 1322 192
rect 1430 188 1434 192
rect 1606 188 1610 192
rect 1630 188 1634 192
rect 1662 188 1666 192
rect 1678 188 1682 192
rect 1790 188 1794 192
rect 1830 188 1834 192
rect 1862 188 1866 192
rect 1942 188 1946 192
rect 2278 188 2282 192
rect 2334 188 2338 192
rect 2382 188 2386 192
rect 2470 188 2474 192
rect 2518 188 2522 192
rect 2566 188 2570 192
rect 2606 188 2610 192
rect 2662 188 2666 192
rect 2694 188 2698 192
rect 2774 188 2778 192
rect 2886 188 2890 192
rect 2942 188 2946 192
rect 3006 188 3010 192
rect 3270 188 3274 192
rect 3414 188 3418 192
rect 3518 188 3522 192
rect 3526 188 3530 192
rect 1206 178 1210 182
rect 1454 178 1458 182
rect 54 168 58 172
rect 294 168 298 172
rect 566 168 570 172
rect 766 168 770 172
rect 862 168 866 172
rect 2374 168 2378 172
rect 2438 168 2442 172
rect 3182 168 3186 172
rect 3398 168 3402 172
rect 310 158 314 162
rect 374 158 378 162
rect 422 158 426 162
rect 454 158 458 162
rect 494 158 498 162
rect 542 158 546 162
rect 598 158 602 162
rect 678 158 682 162
rect 702 158 706 162
rect 6 148 10 152
rect 38 148 42 152
rect 70 148 74 152
rect 134 148 138 152
rect 166 148 170 152
rect 198 148 202 152
rect 222 148 226 152
rect 254 148 258 152
rect 318 148 322 152
rect 358 148 362 152
rect 430 148 434 152
rect 438 148 442 152
rect 510 148 514 152
rect 550 148 554 152
rect 558 148 562 152
rect 582 148 586 152
rect 614 148 618 152
rect 630 148 634 152
rect 646 148 650 152
rect 822 158 826 162
rect 846 158 850 162
rect 878 158 882 162
rect 902 158 906 162
rect 982 158 986 162
rect 1214 158 1218 162
rect 1470 158 1474 162
rect 1550 158 1554 162
rect 1646 158 1650 162
rect 1846 158 1850 162
rect 1878 158 1882 162
rect 1918 158 1922 162
rect 2022 158 2026 162
rect 2046 158 2050 162
rect 2134 158 2138 162
rect 2142 158 2146 162
rect 2262 158 2266 162
rect 2358 158 2362 162
rect 2390 158 2394 162
rect 2454 158 2458 162
rect 2502 158 2506 162
rect 2670 158 2674 162
rect 2758 158 2762 162
rect 2790 158 2794 162
rect 2846 158 2850 162
rect 2902 158 2906 162
rect 2934 158 2938 162
rect 2974 158 2978 162
rect 3030 158 3034 162
rect 3046 158 3050 162
rect 3070 158 3074 162
rect 3118 158 3122 162
rect 3158 158 3162 162
rect 3198 158 3202 162
rect 3206 158 3210 162
rect 3342 158 3346 162
rect 3430 158 3434 162
rect 726 148 730 152
rect 782 148 786 152
rect 806 148 810 152
rect 814 148 818 152
rect 862 148 866 152
rect 950 148 954 152
rect 1054 148 1058 152
rect 1062 148 1066 152
rect 1086 148 1090 152
rect 1102 148 1106 152
rect 1110 148 1114 152
rect 1134 148 1138 152
rect 1150 148 1154 152
rect 1158 148 1162 152
rect 1182 148 1186 152
rect 1262 148 1266 152
rect 1286 148 1290 152
rect 1294 148 1298 152
rect 1310 148 1314 152
rect 1334 148 1338 152
rect 1342 148 1346 152
rect 1350 148 1354 152
rect 1398 148 1402 152
rect 1454 148 1458 152
rect 1478 148 1482 152
rect 1534 148 1538 152
rect 1550 148 1554 152
rect 1606 148 1610 152
rect 1662 148 1666 152
rect 1702 148 1706 152
rect 1726 148 1730 152
rect 1742 148 1746 152
rect 1766 148 1770 152
rect 1830 148 1834 152
rect 1862 148 1866 152
rect 1942 148 1946 152
rect 2038 148 2042 152
rect 2062 148 2066 152
rect 2078 148 2082 152
rect 2118 148 2122 152
rect 2158 148 2162 152
rect 2214 148 2218 152
rect 2222 148 2226 152
rect 2262 148 2266 152
rect 2278 148 2282 152
rect 2302 148 2306 152
rect 2334 148 2338 152
rect 2366 148 2370 152
rect 2398 148 2402 152
rect 2406 148 2410 152
rect 2750 148 2754 152
rect 2774 148 2778 152
rect 2838 148 2842 152
rect 2846 148 2850 152
rect 2862 148 2866 152
rect 2886 148 2890 152
rect 2918 148 2922 152
rect 2926 148 2930 152
rect 2982 148 2986 152
rect 3022 148 3026 152
rect 3030 148 3034 152
rect 3054 148 3058 152
rect 3102 148 3106 152
rect 3126 148 3130 152
rect 3142 148 3146 152
rect 3182 148 3186 152
rect 3246 148 3250 152
rect 3294 148 3298 152
rect 3374 148 3378 152
rect 3422 148 3426 152
rect 3462 148 3466 152
rect 3478 148 3482 152
rect 3550 148 3554 152
rect 30 138 34 142
rect 94 138 98 142
rect 214 138 218 142
rect 286 138 290 142
rect 350 138 354 142
rect 414 138 418 142
rect 446 138 450 142
rect 470 138 474 142
rect 518 138 522 142
rect 526 138 530 142
rect 622 138 626 142
rect 630 138 634 142
rect 662 138 666 142
rect 686 138 690 142
rect 718 138 722 142
rect 734 138 738 142
rect 838 138 842 142
rect 870 138 874 142
rect 894 138 898 142
rect 926 138 930 142
rect 958 138 962 142
rect 998 138 1002 142
rect 1046 138 1050 142
rect 1190 138 1194 142
rect 1246 138 1250 142
rect 1254 138 1258 142
rect 1358 138 1362 142
rect 1382 138 1386 142
rect 1406 138 1410 142
rect 1438 138 1442 142
rect 1446 138 1450 142
rect 1486 138 1490 142
rect 1502 138 1506 142
rect 1526 138 1530 142
rect 1566 138 1570 142
rect 1614 138 1618 142
rect 1670 138 1674 142
rect 1694 138 1698 142
rect 1766 138 1770 142
rect 1814 138 1818 142
rect 1822 138 1826 142
rect 1854 138 1858 142
rect 1886 138 1890 142
rect 1942 138 1946 142
rect 1998 138 2002 142
rect 2006 138 2010 142
rect 2054 138 2058 142
rect 2070 138 2074 142
rect 2086 138 2090 142
rect 2150 138 2154 142
rect 2166 138 2170 142
rect 2190 138 2194 142
rect 2286 138 2290 142
rect 2294 138 2298 142
rect 2414 138 2418 142
rect 2438 138 2442 142
rect 2590 138 2594 142
rect 2646 138 2650 142
rect 2670 138 2674 142
rect 2750 138 2754 142
rect 2782 138 2786 142
rect 2806 138 2810 142
rect 2830 138 2834 142
rect 2870 138 2874 142
rect 2878 138 2882 142
rect 2910 138 2914 142
rect 2950 138 2954 142
rect 2958 138 2962 142
rect 2990 138 2994 142
rect 3014 138 3018 142
rect 3022 138 3026 142
rect 3086 138 3090 142
rect 3110 138 3114 142
rect 3174 138 3178 142
rect 3222 138 3226 142
rect 3326 138 3330 142
rect 3342 138 3346 142
rect 3366 138 3370 142
rect 3422 138 3426 142
rect 3454 138 3458 142
rect 3486 138 3490 142
rect 3510 138 3514 142
rect 3542 138 3546 142
rect 742 128 746 132
rect 766 128 770 132
rect 934 128 938 132
rect 1214 128 1218 132
rect 1238 128 1242 132
rect 1374 128 1378 132
rect 1382 128 1386 132
rect 1398 128 1402 132
rect 1510 128 1514 132
rect 1582 128 1586 132
rect 1638 128 1642 132
rect 1678 128 1682 132
rect 1710 128 1714 132
rect 1910 128 1914 132
rect 1926 128 1930 132
rect 2102 128 2106 132
rect 2134 128 2138 132
rect 2174 128 2178 132
rect 2182 128 2186 132
rect 2206 128 2210 132
rect 2230 128 2234 132
rect 2422 128 2426 132
rect 2478 128 2482 132
rect 2486 128 2490 132
rect 2502 128 2506 132
rect 2590 128 2594 132
rect 2614 128 2618 132
rect 2734 128 2738 132
rect 2814 128 2818 132
rect 2822 128 2826 132
rect 3150 128 3154 132
rect 3158 128 3162 132
rect 3230 128 3234 132
rect 3278 128 3282 132
rect 3318 128 3322 132
rect 3350 128 3354 132
rect 3382 128 3386 132
rect 3462 128 3466 132
rect 3486 128 3490 132
rect 3526 128 3530 132
rect 246 118 250 122
rect 278 118 282 122
rect 390 118 394 122
rect 454 118 458 122
rect 942 118 946 122
rect 1902 118 1906 122
rect 1982 118 1986 122
rect 2454 118 2458 122
rect 2790 118 2794 122
rect 2974 118 2978 122
rect 3206 118 3210 122
rect 3310 118 3314 122
rect 3334 118 3338 122
rect 3430 118 3434 122
rect 190 108 194 112
rect 994 103 998 107
rect 1001 103 1005 107
rect 2026 103 2030 107
rect 2033 103 2037 107
rect 3042 103 3046 107
rect 3049 103 3053 107
rect 150 88 154 92
rect 230 88 234 92
rect 294 88 298 92
rect 326 88 330 92
rect 350 88 354 92
rect 366 88 370 92
rect 422 88 426 92
rect 494 88 498 92
rect 574 88 578 92
rect 622 88 626 92
rect 750 88 754 92
rect 774 88 778 92
rect 790 88 794 92
rect 838 88 842 92
rect 854 88 858 92
rect 886 88 890 92
rect 918 88 922 92
rect 942 88 946 92
rect 1158 88 1162 92
rect 1238 88 1242 92
rect 1462 88 1466 92
rect 1598 88 1602 92
rect 1662 88 1666 92
rect 1726 88 1730 92
rect 1766 88 1770 92
rect 1814 88 1818 92
rect 1870 88 1874 92
rect 1934 88 1938 92
rect 2038 88 2042 92
rect 2094 88 2098 92
rect 2190 88 2194 92
rect 2254 88 2258 92
rect 2270 88 2274 92
rect 2294 88 2298 92
rect 2326 88 2330 92
rect 2350 88 2354 92
rect 2398 88 2402 92
rect 2446 88 2450 92
rect 2510 88 2514 92
rect 2630 88 2634 92
rect 2678 88 2682 92
rect 2742 88 2746 92
rect 2774 88 2778 92
rect 2894 88 2898 92
rect 3006 88 3010 92
rect 3094 88 3098 92
rect 3182 88 3186 92
rect 3222 88 3226 92
rect 3270 88 3274 92
rect 3318 88 3322 92
rect 3358 88 3362 92
rect 54 78 58 82
rect 118 78 122 82
rect 174 79 178 83
rect 374 78 378 82
rect 934 78 938 82
rect 998 78 1002 82
rect 1182 78 1186 82
rect 1214 78 1218 82
rect 1286 78 1290 82
rect 1486 78 1490 82
rect 1494 78 1498 82
rect 1558 78 1562 82
rect 1638 78 1642 82
rect 342 68 346 72
rect 382 68 386 72
rect 398 68 402 72
rect 414 68 418 72
rect 430 68 434 72
rect 462 68 466 72
rect 486 68 490 72
rect 550 68 554 72
rect 582 68 586 72
rect 606 68 610 72
rect 678 68 682 72
rect 726 68 730 72
rect 766 68 770 72
rect 814 68 818 72
rect 822 68 826 72
rect 838 68 842 72
rect 950 68 954 72
rect 966 68 970 72
rect 1030 68 1034 72
rect 1038 68 1042 72
rect 1086 68 1090 72
rect 1102 68 1106 72
rect 1110 68 1114 72
rect 1126 68 1130 72
rect 1174 68 1178 72
rect 1222 68 1226 72
rect 1246 68 1250 72
rect 1294 68 1298 72
rect 1342 68 1346 72
rect 1350 68 1354 72
rect 1366 68 1370 72
rect 1382 68 1386 72
rect 1406 68 1410 72
rect 1438 68 1442 72
rect 1478 68 1482 72
rect 1510 68 1514 72
rect 1542 68 1546 72
rect 1566 68 1570 72
rect 1614 68 1618 72
rect 1654 68 1658 72
rect 1678 78 1682 82
rect 1702 78 1706 82
rect 1694 68 1698 72
rect 1742 78 1746 82
rect 1774 78 1778 82
rect 1878 78 1882 82
rect 1926 78 1930 82
rect 2006 78 2010 82
rect 2022 78 2026 82
rect 1782 68 1786 72
rect 1838 68 1842 72
rect 1846 68 1850 72
rect 1894 68 1898 72
rect 1918 68 1922 72
rect 1942 68 1946 72
rect 1966 68 1970 72
rect 1982 68 1986 72
rect 2030 68 2034 72
rect 2046 68 2050 72
rect 2062 68 2066 72
rect 2110 68 2114 72
rect 2126 68 2130 72
rect 2206 68 2210 72
rect 2286 78 2290 82
rect 2302 78 2306 82
rect 2374 78 2378 82
rect 2406 78 2410 82
rect 2454 78 2458 82
rect 2566 78 2570 82
rect 2686 78 2690 82
rect 2750 78 2754 82
rect 2798 78 2802 82
rect 2942 78 2946 82
rect 3038 78 3042 82
rect 3062 78 3066 82
rect 3134 78 3138 82
rect 3150 78 3154 82
rect 3462 78 3466 82
rect 2238 68 2242 72
rect 2310 68 2314 72
rect 2334 68 2338 72
rect 2390 68 2394 72
rect 2406 68 2410 72
rect 2438 68 2442 72
rect 2478 68 2482 72
rect 2550 68 2554 72
rect 2598 68 2602 72
rect 2654 68 2658 72
rect 2670 68 2674 72
rect 2718 68 2722 72
rect 2726 68 2730 72
rect 2758 68 2762 72
rect 2774 68 2778 72
rect 2798 68 2802 72
rect 2854 68 2858 72
rect 2862 68 2866 72
rect 2910 68 2914 72
rect 2926 68 2930 72
rect 2974 68 2978 72
rect 2982 68 2986 72
rect 3030 68 3034 72
rect 3078 68 3082 72
rect 3126 68 3130 72
rect 3158 68 3162 72
rect 3214 68 3218 72
rect 3230 68 3234 72
rect 3238 68 3242 72
rect 3286 68 3290 72
rect 3342 68 3346 72
rect 3374 68 3378 72
rect 3478 68 3482 72
rect 6 58 10 62
rect 30 58 34 62
rect 38 58 42 62
rect 70 58 74 62
rect 102 58 106 62
rect 134 58 138 62
rect 182 58 186 62
rect 190 58 194 62
rect 214 58 218 62
rect 246 58 250 62
rect 270 58 274 62
rect 310 58 314 62
rect 390 58 394 62
rect 510 58 514 62
rect 534 58 538 62
rect 542 58 546 62
rect 558 58 562 62
rect 638 58 642 62
rect 662 58 666 62
rect 670 58 674 62
rect 718 58 722 62
rect 726 58 730 62
rect 806 58 810 62
rect 870 58 874 62
rect 878 58 882 62
rect 902 58 906 62
rect 958 58 962 62
rect 1022 58 1026 62
rect 1078 58 1082 62
rect 1086 58 1090 62
rect 1222 58 1226 62
rect 1254 58 1258 62
rect 1270 58 1274 62
rect 1326 58 1330 62
rect 1358 58 1362 62
rect 1414 58 1418 62
rect 1430 58 1434 62
rect 1446 58 1450 62
rect 1470 58 1474 62
rect 1518 58 1522 62
rect 1534 58 1538 62
rect 1622 58 1626 62
rect 1798 58 1802 62
rect 1854 58 1858 62
rect 1910 58 1914 62
rect 1950 58 1954 62
rect 1974 58 1978 62
rect 1990 58 1994 62
rect 2054 58 2058 62
rect 2150 58 2154 62
rect 2158 58 2162 62
rect 2222 58 2226 62
rect 2230 58 2234 62
rect 2262 58 2266 62
rect 2286 58 2290 62
rect 2358 58 2362 62
rect 2382 58 2386 62
rect 2430 58 2434 62
rect 2470 58 2474 62
rect 2550 58 2554 62
rect 2598 58 2602 62
rect 2606 58 2610 62
rect 2646 58 2650 62
rect 2662 58 2666 62
rect 2694 58 2698 62
rect 2710 58 2714 62
rect 2726 58 2730 62
rect 2782 58 2786 62
rect 2918 58 2922 62
rect 2950 58 2954 62
rect 2966 58 2970 62
rect 3134 58 3138 62
rect 3294 58 3298 62
rect 3334 58 3338 62
rect 3381 58 3385 62
rect 3526 58 3530 62
rect 262 48 266 52
rect 358 48 362 52
rect 406 48 410 52
rect 430 48 434 52
rect 454 48 458 52
rect 478 48 482 52
rect 598 48 602 52
rect 622 48 626 52
rect 646 48 650 52
rect 694 48 698 52
rect 782 48 786 52
rect 790 48 794 52
rect 838 48 842 52
rect 862 48 866 52
rect 982 48 986 52
rect 1054 48 1058 52
rect 1118 48 1122 52
rect 1238 48 1242 52
rect 1254 48 1258 52
rect 1270 48 1274 52
rect 1374 48 1378 52
rect 1398 48 1402 52
rect 1430 48 1434 52
rect 1462 48 1466 52
rect 1806 48 1810 52
rect 1822 48 1826 52
rect 1870 48 1874 52
rect 1958 48 1962 52
rect 2118 48 2122 52
rect 2254 48 2258 52
rect 2326 48 2330 52
rect 2414 48 2418 52
rect 2590 48 2594 52
rect 2622 48 2626 52
rect 2774 48 2778 52
rect 2950 48 2954 52
rect 3214 48 3218 52
rect 3318 48 3322 52
rect 3526 48 3530 52
rect 86 38 90 42
rect 702 38 706 42
rect 1078 38 1082 42
rect 1838 38 1842 42
rect 2838 38 2842 42
rect 2966 38 2970 42
rect 3310 38 3314 42
rect 446 28 450 32
rect 718 28 722 32
rect 2366 28 2370 32
rect 2606 28 2610 32
rect 166 18 170 22
rect 206 18 210 22
rect 1558 18 1562 22
rect 2134 18 2138 22
rect 3526 18 3530 22
rect 482 3 486 7
rect 489 3 493 7
rect 1514 3 1518 7
rect 1521 3 1525 7
rect 2538 3 2542 7
rect 2545 3 2549 7
<< metal2 >>
rect 190 3331 194 3332
rect 334 3331 338 3332
rect 182 3328 194 3331
rect 326 3328 338 3331
rect 406 3331 410 3332
rect 406 3328 417 3331
rect 182 3292 185 3328
rect 326 3292 329 3328
rect 414 3292 417 3328
rect 502 3328 506 3332
rect 526 3331 530 3332
rect 526 3328 537 3331
rect 502 3292 505 3328
rect 534 3292 537 3328
rect 606 3328 610 3332
rect 630 3328 634 3332
rect 646 3328 650 3332
rect 670 3328 674 3332
rect 694 3328 698 3332
rect 710 3328 714 3332
rect 734 3328 738 3332
rect 750 3328 754 3332
rect 854 3328 858 3332
rect 1022 3328 1026 3332
rect 1054 3328 1058 3332
rect 1142 3328 1146 3332
rect 1230 3328 1234 3332
rect 1246 3328 1250 3332
rect 1286 3328 1290 3332
rect 1350 3328 1354 3332
rect 1374 3328 1378 3332
rect 1390 3328 1394 3332
rect 1414 3328 1418 3332
rect 1430 3328 1434 3332
rect 1534 3328 1538 3332
rect 1550 3328 1554 3332
rect 1574 3328 1578 3332
rect 1598 3328 1602 3332
rect 1646 3328 1650 3332
rect 1670 3328 1674 3332
rect 1686 3331 1690 3332
rect 1678 3328 1690 3331
rect 1702 3328 1706 3332
rect 1726 3328 1730 3332
rect 1742 3328 1746 3332
rect 1854 3331 1858 3332
rect 1854 3328 1865 3331
rect 606 3302 609 3328
rect 630 3292 633 3328
rect 110 3272 113 3278
rect 94 3263 97 3268
rect 6 3242 9 3248
rect 30 3242 33 3248
rect 126 3222 129 3258
rect 134 3222 137 3268
rect 142 3262 145 3268
rect 158 3252 161 3258
rect 174 3232 177 3278
rect 198 3262 201 3268
rect 222 3262 225 3278
rect 254 3272 257 3278
rect 206 3252 209 3258
rect 214 3242 217 3248
rect 102 3192 105 3218
rect 174 3192 177 3218
rect 90 3168 94 3171
rect 78 3162 81 3168
rect 34 3158 38 3161
rect 114 3158 118 3161
rect 18 3148 25 3151
rect 10 3138 14 3141
rect 22 3132 25 3148
rect 30 3142 33 3148
rect 38 3142 41 3148
rect 22 3082 25 3128
rect 38 3082 41 3138
rect 46 3092 49 3158
rect 98 3148 102 3151
rect 134 3142 137 3148
rect 150 3142 153 3148
rect 82 3138 86 3141
rect 166 3138 174 3141
rect 54 3122 57 3128
rect 78 3092 81 3138
rect 158 3132 161 3138
rect 118 3122 121 3128
rect 142 3122 145 3128
rect 166 3122 169 3138
rect 174 3122 177 3128
rect 166 3092 169 3118
rect 6 3072 9 3078
rect 54 3072 57 3088
rect 134 3082 137 3088
rect 34 3068 38 3071
rect 6 3052 9 3068
rect 62 3062 65 3078
rect 74 3068 78 3071
rect 26 3058 30 3061
rect 22 2962 25 3018
rect 38 2952 41 3018
rect 46 2942 49 3018
rect 78 2952 81 3048
rect 86 3042 89 3078
rect 142 3062 145 3068
rect 102 2972 105 3058
rect 118 3042 121 3058
rect 134 2962 137 2968
rect 86 2952 89 2958
rect 58 2948 62 2951
rect 42 2938 46 2941
rect 90 2938 94 2941
rect 58 2928 62 2931
rect 106 2928 110 2931
rect 6 2911 9 2928
rect 18 2918 22 2921
rect 6 2908 17 2911
rect 14 2892 17 2908
rect 6 2852 9 2878
rect 22 2872 25 2878
rect 38 2862 41 2928
rect 54 2892 57 2918
rect 70 2892 73 2918
rect 78 2892 81 2928
rect 118 2921 121 2928
rect 110 2918 121 2921
rect 134 2922 137 2948
rect 142 2932 145 3058
rect 150 2952 153 3058
rect 174 2992 177 3068
rect 182 2962 185 3148
rect 202 3138 206 3141
rect 206 3072 209 3128
rect 222 3122 225 3258
rect 254 3152 257 3268
rect 266 3258 270 3261
rect 318 3222 321 3268
rect 346 3258 350 3261
rect 390 3261 393 3278
rect 458 3268 462 3271
rect 390 3258 398 3261
rect 318 3172 321 3218
rect 314 3148 318 3151
rect 278 3132 281 3147
rect 294 3142 297 3148
rect 218 3118 222 3121
rect 294 3092 297 3128
rect 238 3072 241 3078
rect 286 3072 289 3088
rect 194 3068 198 3071
rect 198 3062 201 3068
rect 210 3058 214 3061
rect 222 3052 225 3068
rect 246 3062 249 3068
rect 310 3062 313 3118
rect 318 3082 321 3138
rect 326 3132 329 3228
rect 334 3192 337 3258
rect 346 3248 350 3251
rect 358 3242 361 3248
rect 366 3192 369 3258
rect 398 3192 401 3258
rect 422 3252 425 3258
rect 430 3252 433 3258
rect 470 3242 473 3278
rect 478 3262 481 3268
rect 606 3263 609 3268
rect 518 3242 521 3258
rect 622 3252 625 3268
rect 638 3242 641 3258
rect 546 3238 550 3241
rect 326 3082 329 3128
rect 334 3062 337 3158
rect 342 3152 345 3168
rect 398 3148 406 3151
rect 362 3128 366 3131
rect 354 3088 358 3091
rect 342 3062 345 3068
rect 254 3052 257 3058
rect 334 3052 337 3058
rect 194 3048 198 3051
rect 270 3042 273 3048
rect 206 3032 209 3038
rect 238 3032 241 3038
rect 190 2952 193 2958
rect 154 2948 158 2951
rect 206 2942 209 3028
rect 286 2992 289 3048
rect 350 2992 353 3078
rect 358 3042 361 3078
rect 366 3062 369 3118
rect 382 3082 385 3128
rect 398 3092 401 3148
rect 410 3138 414 3141
rect 446 3122 449 3138
rect 462 3132 465 3218
rect 480 3203 482 3207
rect 486 3203 489 3207
rect 493 3203 496 3207
rect 494 3152 497 3188
rect 546 3148 550 3151
rect 470 3082 473 3118
rect 494 3092 497 3148
rect 502 3132 505 3148
rect 522 3138 526 3141
rect 478 3072 481 3078
rect 274 2958 278 2961
rect 370 2958 374 2961
rect 234 2948 238 2951
rect 254 2942 257 2958
rect 266 2948 270 2951
rect 170 2928 174 2931
rect 70 2862 73 2878
rect 86 2872 89 2878
rect 94 2872 97 2878
rect 70 2852 73 2858
rect 102 2852 105 2918
rect 110 2902 113 2918
rect 142 2912 145 2928
rect 150 2912 153 2918
rect 110 2882 113 2898
rect 182 2881 185 2938
rect 202 2928 206 2931
rect 190 2892 193 2928
rect 198 2882 201 2918
rect 214 2902 217 2928
rect 230 2922 233 2938
rect 230 2882 233 2918
rect 238 2882 241 2908
rect 246 2882 249 2918
rect 182 2878 190 2881
rect 158 2872 161 2878
rect 146 2868 150 2871
rect 110 2862 113 2868
rect 174 2862 177 2868
rect 114 2848 118 2851
rect 6 2742 9 2848
rect 14 2792 17 2848
rect 134 2832 137 2858
rect 150 2842 153 2848
rect 30 2792 33 2808
rect 94 2792 97 2828
rect 118 2792 121 2818
rect 134 2772 137 2818
rect 166 2812 169 2858
rect 38 2758 46 2761
rect 82 2758 86 2761
rect 162 2758 166 2761
rect 190 2761 193 2878
rect 234 2868 238 2871
rect 262 2862 265 2898
rect 278 2892 281 2898
rect 286 2882 289 2958
rect 390 2952 393 2958
rect 370 2948 374 2951
rect 310 2942 313 2948
rect 342 2942 345 2948
rect 350 2942 353 2948
rect 338 2938 342 2941
rect 386 2938 390 2941
rect 294 2912 297 2938
rect 294 2882 297 2888
rect 302 2882 305 2898
rect 210 2858 214 2861
rect 250 2858 254 2861
rect 202 2848 206 2851
rect 274 2848 278 2851
rect 286 2832 289 2878
rect 302 2842 305 2848
rect 190 2758 198 2761
rect 274 2758 278 2761
rect 10 2738 14 2741
rect 22 2732 25 2738
rect 6 2682 9 2698
rect 14 2682 17 2718
rect 30 2702 33 2748
rect 38 2672 41 2758
rect 58 2748 62 2751
rect 146 2748 150 2751
rect 162 2748 166 2751
rect 154 2738 158 2741
rect 54 2732 57 2738
rect 134 2732 137 2738
rect 54 2681 57 2728
rect 94 2682 97 2688
rect 54 2678 62 2681
rect 26 2668 30 2671
rect 54 2662 57 2678
rect 78 2672 81 2678
rect 62 2662 65 2668
rect 10 2658 14 2661
rect 26 2658 30 2661
rect 90 2658 94 2661
rect 30 2652 33 2658
rect 6 2562 9 2608
rect 14 2592 17 2618
rect 6 2542 9 2558
rect 30 2542 33 2628
rect 38 2592 41 2658
rect 46 2542 49 2658
rect 78 2652 81 2658
rect 94 2612 97 2658
rect 102 2632 105 2678
rect 118 2662 121 2698
rect 158 2672 161 2678
rect 174 2672 177 2758
rect 302 2752 305 2758
rect 310 2752 313 2938
rect 398 2932 401 3068
rect 462 3062 465 3068
rect 442 3058 446 3061
rect 414 2982 417 3058
rect 426 3048 430 3051
rect 454 3032 457 3058
rect 462 2992 465 3058
rect 470 3052 473 3058
rect 542 3052 545 3138
rect 558 3122 561 3238
rect 582 3162 585 3168
rect 638 3162 641 3168
rect 570 3158 574 3161
rect 602 3158 606 3161
rect 602 3148 606 3151
rect 634 3148 638 3151
rect 582 3142 585 3148
rect 570 3138 574 3141
rect 574 3122 577 3138
rect 558 3072 561 3118
rect 566 3102 569 3118
rect 598 3112 601 3148
rect 606 3132 609 3138
rect 610 3088 614 3091
rect 598 3082 601 3088
rect 622 3082 625 3128
rect 646 3112 649 3328
rect 670 3302 673 3328
rect 694 3302 697 3328
rect 654 3222 657 3278
rect 690 3268 694 3271
rect 666 3258 670 3261
rect 678 3212 681 3268
rect 702 3262 705 3298
rect 710 3272 713 3328
rect 734 3302 737 3328
rect 690 3258 694 3261
rect 670 3152 673 3158
rect 682 3148 689 3151
rect 658 3138 662 3141
rect 646 3072 649 3108
rect 606 3068 614 3071
rect 562 3059 566 3062
rect 480 3003 482 3007
rect 486 3003 489 3007
rect 493 3003 496 3007
rect 518 2992 521 3018
rect 434 2948 438 2951
rect 538 2948 542 2951
rect 406 2942 409 2948
rect 338 2928 342 2931
rect 434 2928 438 2931
rect 318 2872 321 2878
rect 326 2872 329 2918
rect 406 2902 409 2928
rect 346 2888 350 2891
rect 334 2862 337 2868
rect 350 2852 353 2868
rect 374 2862 377 2868
rect 362 2848 366 2851
rect 326 2792 329 2848
rect 374 2802 377 2818
rect 382 2792 385 2868
rect 414 2862 417 2918
rect 446 2912 449 2948
rect 470 2942 473 2948
rect 558 2942 561 2948
rect 454 2902 457 2928
rect 478 2912 481 2928
rect 426 2878 430 2881
rect 450 2878 454 2881
rect 462 2872 465 2888
rect 470 2882 473 2888
rect 426 2868 430 2871
rect 394 2858 398 2861
rect 410 2848 414 2851
rect 406 2792 409 2828
rect 250 2748 254 2751
rect 282 2748 286 2751
rect 330 2748 334 2751
rect 342 2748 350 2751
rect 378 2748 382 2751
rect 186 2738 190 2741
rect 190 2712 193 2718
rect 198 2702 201 2748
rect 270 2742 273 2748
rect 314 2738 326 2741
rect 206 2732 209 2738
rect 222 2732 225 2738
rect 278 2732 281 2738
rect 230 2721 233 2728
rect 222 2718 233 2721
rect 198 2692 201 2698
rect 222 2692 225 2718
rect 214 2682 217 2688
rect 190 2672 193 2678
rect 206 2672 209 2678
rect 154 2668 158 2671
rect 118 2642 121 2648
rect 126 2632 129 2668
rect 166 2662 169 2668
rect 206 2662 209 2668
rect 150 2652 153 2658
rect 166 2652 169 2658
rect 186 2648 190 2651
rect 102 2592 105 2598
rect 134 2572 137 2618
rect 174 2582 177 2588
rect 58 2558 62 2561
rect 78 2552 81 2568
rect 126 2562 129 2568
rect 30 2522 33 2538
rect 70 2532 73 2538
rect 78 2532 81 2548
rect 110 2532 113 2548
rect 134 2532 137 2548
rect 182 2542 185 2618
rect 214 2582 217 2678
rect 222 2652 225 2688
rect 250 2678 254 2681
rect 230 2662 233 2678
rect 262 2662 265 2678
rect 270 2672 273 2698
rect 278 2692 281 2718
rect 294 2702 297 2738
rect 326 2702 329 2728
rect 342 2712 345 2748
rect 362 2738 369 2741
rect 358 2732 361 2738
rect 350 2722 353 2728
rect 366 2722 369 2738
rect 286 2672 289 2678
rect 318 2672 321 2698
rect 390 2691 393 2778
rect 398 2732 401 2768
rect 446 2762 449 2858
rect 454 2852 457 2858
rect 462 2752 465 2848
rect 478 2832 481 2858
rect 490 2848 494 2851
rect 480 2803 482 2807
rect 486 2803 489 2807
rect 493 2803 496 2807
rect 458 2748 462 2751
rect 490 2748 494 2751
rect 438 2742 441 2748
rect 502 2742 505 2938
rect 558 2921 561 2938
rect 582 2932 585 3068
rect 590 2942 593 3028
rect 570 2928 574 2931
rect 598 2931 601 3058
rect 606 3042 609 3068
rect 670 3062 673 3118
rect 678 3082 681 3128
rect 686 3122 689 3148
rect 702 3142 705 3258
rect 726 3252 729 3278
rect 734 3262 737 3268
rect 742 3262 745 3268
rect 742 3242 745 3258
rect 750 3232 753 3328
rect 774 3282 777 3288
rect 782 3282 785 3288
rect 854 3272 857 3328
rect 992 3303 994 3307
rect 998 3303 1001 3307
rect 1005 3303 1008 3307
rect 1022 3302 1025 3328
rect 1054 3302 1057 3328
rect 1142 3302 1145 3328
rect 1230 3302 1233 3328
rect 930 3288 934 3291
rect 1018 3288 1025 3291
rect 894 3282 897 3288
rect 1022 3282 1025 3288
rect 882 3278 886 3281
rect 898 3278 902 3281
rect 962 3278 966 3281
rect 1178 3278 1182 3281
rect 770 3268 774 3271
rect 858 3268 862 3271
rect 762 3258 766 3261
rect 790 3252 793 3258
rect 710 3172 713 3178
rect 718 3162 721 3218
rect 734 3142 737 3168
rect 790 3162 793 3248
rect 818 3168 822 3171
rect 798 3162 801 3168
rect 830 3162 833 3168
rect 742 3152 745 3158
rect 838 3152 841 3178
rect 862 3152 865 3258
rect 870 3242 873 3268
rect 886 3262 889 3268
rect 910 3262 913 3268
rect 958 3262 961 3268
rect 922 3258 926 3261
rect 902 3251 905 3258
rect 942 3252 945 3258
rect 902 3248 926 3251
rect 910 3192 913 3208
rect 934 3192 937 3238
rect 810 3148 814 3151
rect 834 3148 838 3151
rect 766 3142 769 3148
rect 774 3142 777 3148
rect 798 3142 801 3148
rect 862 3142 865 3148
rect 778 3138 782 3141
rect 698 3128 702 3131
rect 762 3128 766 3131
rect 718 3122 721 3128
rect 726 3122 729 3128
rect 718 3082 721 3118
rect 750 3112 753 3128
rect 678 3072 681 3078
rect 618 3058 622 3061
rect 626 3048 630 3051
rect 686 3032 689 3068
rect 670 3002 673 3018
rect 670 2962 673 2968
rect 634 2948 638 2951
rect 622 2942 625 2948
rect 610 2938 614 2941
rect 630 2932 633 2938
rect 590 2928 601 2931
rect 610 2928 614 2931
rect 558 2918 569 2921
rect 566 2892 569 2918
rect 574 2891 577 2918
rect 590 2892 593 2928
rect 574 2888 585 2891
rect 550 2872 553 2878
rect 514 2858 518 2861
rect 510 2752 513 2818
rect 542 2812 545 2858
rect 558 2802 561 2878
rect 574 2872 577 2878
rect 582 2871 585 2888
rect 582 2868 593 2871
rect 582 2842 585 2858
rect 590 2852 593 2868
rect 598 2862 601 2918
rect 614 2852 617 2868
rect 590 2792 593 2798
rect 554 2748 558 2751
rect 382 2688 393 2691
rect 326 2662 329 2668
rect 222 2592 225 2638
rect 230 2592 233 2658
rect 238 2612 241 2658
rect 294 2652 297 2658
rect 262 2592 265 2608
rect 190 2552 193 2568
rect 242 2558 246 2561
rect 162 2538 166 2541
rect 42 2528 46 2531
rect 6 2492 9 2508
rect 14 2482 17 2518
rect 54 2502 57 2518
rect 10 2468 14 2471
rect 18 2458 22 2461
rect 6 2362 9 2398
rect 6 2252 9 2318
rect 14 2172 17 2418
rect 30 2382 33 2478
rect 38 2462 41 2498
rect 70 2492 73 2518
rect 46 2482 49 2488
rect 54 2472 57 2478
rect 38 2372 41 2458
rect 54 2452 57 2468
rect 62 2432 65 2468
rect 54 2362 57 2368
rect 62 2362 65 2368
rect 34 2348 38 2351
rect 34 2338 38 2341
rect 22 2262 25 2338
rect 30 2272 33 2338
rect 46 2292 49 2358
rect 78 2352 81 2468
rect 78 2332 81 2348
rect 86 2342 89 2518
rect 94 2472 97 2528
rect 110 2522 113 2528
rect 158 2522 161 2528
rect 150 2512 153 2518
rect 142 2482 145 2508
rect 158 2492 161 2498
rect 134 2472 137 2478
rect 126 2462 129 2468
rect 94 2442 97 2448
rect 94 2342 97 2378
rect 102 2362 105 2458
rect 110 2432 113 2458
rect 122 2448 126 2451
rect 134 2442 137 2468
rect 142 2462 145 2478
rect 150 2472 153 2478
rect 166 2462 169 2518
rect 174 2482 177 2518
rect 198 2492 201 2508
rect 206 2502 209 2518
rect 214 2491 217 2538
rect 222 2522 225 2548
rect 262 2502 265 2548
rect 270 2542 273 2628
rect 310 2622 313 2658
rect 302 2552 305 2578
rect 318 2562 321 2658
rect 334 2582 337 2658
rect 278 2542 281 2548
rect 326 2542 329 2568
rect 290 2538 294 2541
rect 270 2512 273 2538
rect 210 2488 217 2491
rect 222 2492 225 2498
rect 182 2472 185 2488
rect 206 2482 209 2488
rect 190 2462 193 2468
rect 170 2458 174 2461
rect 154 2448 158 2451
rect 118 2362 121 2368
rect 114 2358 118 2361
rect 126 2352 129 2358
rect 134 2352 137 2428
rect 158 2352 161 2438
rect 174 2362 177 2368
rect 102 2342 105 2348
rect 54 2272 57 2318
rect 62 2302 65 2318
rect 94 2281 97 2338
rect 86 2278 97 2281
rect 102 2282 105 2298
rect 118 2281 121 2318
rect 126 2281 129 2288
rect 118 2278 129 2281
rect 86 2272 89 2278
rect 38 2262 41 2268
rect 94 2262 97 2268
rect 102 2262 105 2278
rect 30 2252 33 2258
rect 94 2252 97 2258
rect 10 2148 14 2151
rect 22 2132 25 2218
rect 30 2152 33 2158
rect 54 2152 57 2238
rect 78 2202 81 2218
rect 110 2182 113 2218
rect 118 2171 121 2268
rect 126 2262 129 2278
rect 134 2272 137 2348
rect 150 2312 153 2318
rect 150 2262 153 2288
rect 174 2262 177 2318
rect 182 2272 185 2338
rect 190 2332 193 2348
rect 198 2342 201 2478
rect 210 2458 214 2461
rect 230 2442 233 2478
rect 238 2442 241 2448
rect 254 2432 257 2468
rect 278 2462 281 2528
rect 286 2522 289 2528
rect 334 2522 337 2548
rect 350 2542 353 2678
rect 374 2662 377 2678
rect 382 2662 385 2688
rect 390 2672 393 2678
rect 406 2672 409 2688
rect 414 2682 417 2738
rect 482 2728 486 2731
rect 422 2711 425 2728
rect 434 2718 441 2721
rect 422 2708 433 2711
rect 430 2692 433 2708
rect 414 2662 417 2668
rect 358 2582 361 2598
rect 358 2552 361 2578
rect 390 2572 393 2618
rect 398 2592 401 2598
rect 406 2551 409 2638
rect 422 2612 425 2668
rect 438 2662 441 2718
rect 470 2712 473 2718
rect 510 2712 513 2738
rect 534 2732 537 2738
rect 510 2682 513 2698
rect 518 2692 521 2698
rect 526 2682 529 2728
rect 450 2678 457 2681
rect 462 2662 465 2678
rect 442 2648 446 2651
rect 450 2648 457 2651
rect 446 2552 449 2568
rect 454 2562 457 2648
rect 462 2632 465 2658
rect 478 2642 481 2648
rect 480 2603 482 2607
rect 486 2603 489 2607
rect 493 2603 496 2607
rect 510 2582 513 2678
rect 526 2672 529 2678
rect 510 2552 513 2558
rect 402 2548 409 2551
rect 426 2548 430 2551
rect 374 2542 377 2548
rect 322 2518 326 2521
rect 286 2472 289 2518
rect 302 2472 305 2508
rect 342 2482 345 2498
rect 294 2462 297 2468
rect 326 2462 329 2478
rect 282 2458 286 2461
rect 238 2362 241 2378
rect 214 2352 217 2358
rect 222 2322 225 2338
rect 230 2322 233 2358
rect 198 2262 201 2318
rect 222 2262 225 2298
rect 134 2252 137 2258
rect 182 2252 185 2258
rect 230 2252 233 2258
rect 110 2168 121 2171
rect 110 2162 113 2168
rect 150 2162 153 2218
rect 166 2212 169 2218
rect 190 2162 193 2168
rect 194 2158 198 2161
rect 70 2152 73 2158
rect 118 2152 121 2158
rect 206 2152 209 2218
rect 230 2192 233 2248
rect 214 2162 217 2178
rect 90 2148 94 2151
rect 10 2128 14 2131
rect 6 2042 9 2068
rect 18 2048 22 2051
rect 6 1942 9 2038
rect 14 1952 17 2048
rect 38 1952 41 2118
rect 50 2068 54 2071
rect 46 2042 49 2058
rect 62 2052 65 2148
rect 70 2072 73 2148
rect 82 2138 86 2141
rect 162 2138 166 2141
rect 178 2138 182 2141
rect 94 2132 97 2138
rect 86 2072 89 2078
rect 78 2052 81 2058
rect 94 2052 97 2058
rect 110 2052 113 2118
rect 118 2032 121 2118
rect 126 2082 129 2108
rect 134 2052 137 2088
rect 150 2062 153 2138
rect 198 2132 201 2138
rect 162 2128 169 2131
rect 158 2072 161 2118
rect 166 2092 169 2128
rect 166 2072 169 2078
rect 174 2062 177 2128
rect 34 1938 38 1941
rect 6 1872 9 1938
rect 6 1732 9 1758
rect 6 1662 9 1718
rect 14 1581 17 1878
rect 30 1872 33 1918
rect 46 1881 49 2018
rect 70 1972 73 2018
rect 70 1932 73 1958
rect 38 1878 49 1881
rect 30 1852 33 1858
rect 38 1762 41 1878
rect 78 1871 81 2028
rect 94 1992 97 2018
rect 94 1962 97 1988
rect 118 1972 121 2018
rect 90 1948 94 1951
rect 130 1948 134 1951
rect 70 1868 81 1871
rect 98 1938 102 1941
rect 122 1938 126 1941
rect 86 1872 89 1938
rect 94 1882 97 1898
rect 102 1882 105 1888
rect 46 1862 49 1868
rect 70 1862 73 1868
rect 62 1812 65 1818
rect 70 1802 73 1858
rect 78 1842 81 1858
rect 98 1848 102 1851
rect 62 1762 65 1768
rect 22 1742 25 1748
rect 30 1742 33 1758
rect 38 1752 41 1758
rect 58 1738 62 1741
rect 38 1732 41 1738
rect 30 1692 33 1708
rect 38 1662 41 1668
rect 6 1578 17 1581
rect 6 1482 9 1578
rect 14 1562 17 1568
rect 34 1548 38 1551
rect 46 1551 49 1658
rect 62 1651 65 1718
rect 70 1662 73 1768
rect 78 1752 81 1838
rect 86 1762 89 1818
rect 110 1782 113 1918
rect 118 1862 121 1908
rect 142 1902 145 2058
rect 150 2042 153 2058
rect 174 2032 177 2058
rect 190 2052 193 2118
rect 198 2062 201 2068
rect 206 2051 209 2118
rect 202 2048 209 2051
rect 214 2062 217 2128
rect 238 2092 241 2318
rect 246 2262 249 2278
rect 254 2252 257 2348
rect 270 2262 273 2458
rect 318 2442 321 2448
rect 350 2412 353 2518
rect 366 2462 369 2538
rect 382 2532 385 2548
rect 374 2522 377 2528
rect 398 2472 401 2548
rect 470 2542 473 2548
rect 518 2542 521 2608
rect 526 2552 529 2658
rect 534 2652 537 2658
rect 534 2592 537 2648
rect 526 2542 529 2548
rect 534 2542 537 2548
rect 542 2542 545 2748
rect 550 2692 553 2708
rect 558 2702 561 2738
rect 566 2732 569 2748
rect 582 2742 585 2748
rect 598 2742 601 2848
rect 622 2842 625 2848
rect 618 2788 622 2791
rect 610 2738 614 2741
rect 562 2698 569 2701
rect 558 2672 561 2678
rect 566 2662 569 2698
rect 582 2662 585 2728
rect 590 2672 593 2688
rect 598 2662 601 2738
rect 622 2732 625 2768
rect 630 2742 633 2928
rect 646 2872 649 2908
rect 654 2902 657 2918
rect 670 2882 673 2948
rect 678 2932 681 2938
rect 686 2932 689 2958
rect 694 2952 697 3058
rect 710 2962 713 3008
rect 718 2982 721 3038
rect 734 3022 737 3078
rect 754 3058 758 3061
rect 774 3052 777 3098
rect 726 2992 729 3018
rect 734 3012 737 3018
rect 686 2892 689 2928
rect 694 2922 697 2938
rect 702 2931 705 2948
rect 710 2942 713 2958
rect 726 2952 729 2958
rect 734 2942 737 2998
rect 742 2952 745 3018
rect 766 2962 769 3018
rect 782 2992 785 3048
rect 790 3031 793 3138
rect 806 3132 809 3138
rect 850 3128 854 3131
rect 846 3102 849 3118
rect 814 3082 817 3098
rect 826 3088 830 3091
rect 802 3058 806 3061
rect 798 3042 801 3048
rect 830 3032 833 3068
rect 846 3062 849 3078
rect 790 3028 801 3031
rect 786 2958 790 2961
rect 702 2928 713 2931
rect 710 2882 713 2928
rect 718 2922 721 2928
rect 750 2892 753 2938
rect 790 2932 793 2938
rect 762 2918 766 2921
rect 774 2882 777 2928
rect 798 2892 801 3028
rect 822 2942 825 2948
rect 810 2938 814 2941
rect 830 2941 833 2998
rect 838 2962 841 3058
rect 846 2962 849 3058
rect 854 2972 857 3128
rect 862 3102 865 3128
rect 862 3082 865 3098
rect 878 3091 881 3158
rect 898 3138 905 3141
rect 874 3088 881 3091
rect 902 3092 905 3138
rect 910 3112 913 3128
rect 918 3122 921 3158
rect 950 3152 953 3158
rect 958 3152 961 3258
rect 966 3172 969 3218
rect 974 3192 977 3258
rect 998 3182 1001 3278
rect 1006 3262 1009 3268
rect 1014 3192 1017 3278
rect 1038 3262 1041 3268
rect 1078 3262 1081 3268
rect 1086 3262 1089 3278
rect 1050 3258 1054 3261
rect 1070 3252 1073 3258
rect 1022 3242 1025 3248
rect 1054 3242 1057 3248
rect 1070 3232 1073 3238
rect 1078 3202 1081 3258
rect 1094 3232 1097 3268
rect 1106 3258 1110 3261
rect 1118 3252 1121 3278
rect 1246 3262 1249 3328
rect 1286 3302 1289 3328
rect 1350 3302 1353 3328
rect 1354 3288 1358 3291
rect 1270 3262 1273 3288
rect 1194 3258 1198 3261
rect 1330 3258 1334 3261
rect 1294 3242 1297 3258
rect 1326 3242 1329 3248
rect 1110 3192 1113 3198
rect 1190 3162 1193 3168
rect 942 3122 945 3138
rect 966 3132 969 3138
rect 974 3122 977 3148
rect 1022 3142 1025 3158
rect 1114 3148 1118 3151
rect 990 3132 993 3138
rect 1038 3122 1041 3147
rect 918 3102 921 3118
rect 870 3082 873 3088
rect 922 3078 926 3081
rect 886 2972 889 3058
rect 910 3012 913 3078
rect 918 3052 921 3058
rect 918 2992 921 3048
rect 934 3022 937 3068
rect 950 3061 953 3118
rect 992 3103 994 3107
rect 998 3103 1001 3107
rect 1005 3103 1008 3107
rect 946 3058 953 3061
rect 958 3082 961 3088
rect 958 3062 961 3078
rect 966 3072 969 3098
rect 1026 3058 1030 3061
rect 950 3042 953 3048
rect 966 2992 969 3058
rect 1038 3052 1041 3068
rect 1046 3022 1049 3068
rect 1054 3062 1057 3148
rect 1062 3142 1065 3148
rect 1158 3142 1161 3148
rect 1166 3142 1169 3148
rect 1130 3138 1134 3141
rect 1062 3092 1065 3138
rect 1070 3072 1073 3128
rect 1118 3122 1121 3128
rect 1098 3118 1102 3121
rect 1138 3118 1142 3121
rect 1150 3082 1153 3128
rect 1182 3122 1185 3158
rect 1198 3151 1201 3228
rect 1262 3192 1265 3198
rect 1250 3168 1254 3171
rect 1206 3162 1209 3168
rect 1238 3152 1241 3158
rect 1198 3148 1209 3151
rect 1250 3148 1254 3151
rect 1190 3142 1193 3148
rect 1206 3092 1209 3148
rect 1270 3142 1273 3178
rect 1342 3172 1345 3268
rect 1374 3262 1377 3328
rect 1286 3152 1289 3158
rect 1310 3152 1313 3158
rect 1358 3152 1361 3258
rect 1366 3252 1369 3258
rect 1382 3222 1385 3278
rect 1354 3148 1358 3151
rect 1278 3142 1281 3148
rect 1342 3142 1345 3148
rect 1374 3142 1377 3148
rect 1382 3142 1385 3158
rect 1214 3132 1217 3138
rect 1230 3102 1233 3128
rect 1230 3092 1233 3098
rect 1158 3082 1161 3088
rect 1146 3078 1150 3081
rect 1210 3078 1214 3081
rect 1078 3072 1081 3078
rect 1102 3072 1105 3078
rect 1134 3072 1137 3078
rect 1142 3068 1150 3071
rect 1058 3058 1062 3061
rect 1078 3042 1081 3068
rect 1142 3062 1145 3068
rect 1122 3058 1126 3061
rect 1154 3058 1190 3061
rect 1122 3048 1126 3051
rect 1086 3042 1089 3048
rect 1094 3022 1097 3048
rect 1222 3042 1225 3078
rect 1238 3072 1241 3128
rect 1294 3112 1297 3138
rect 1254 3082 1257 3098
rect 1286 3072 1289 3078
rect 1326 3072 1329 3088
rect 1350 3082 1353 3128
rect 1366 3112 1369 3128
rect 1390 3082 1393 3328
rect 1414 3302 1417 3328
rect 1430 3242 1433 3328
rect 1454 3262 1457 3268
rect 1398 3232 1401 3238
rect 1398 3182 1401 3228
rect 1402 3168 1406 3171
rect 1430 3152 1433 3208
rect 1462 3192 1465 3278
rect 1478 3262 1481 3268
rect 1486 3262 1489 3268
rect 1506 3258 1510 3261
rect 1470 3252 1473 3258
rect 1478 3212 1481 3258
rect 1490 3248 1494 3251
rect 1510 3242 1513 3248
rect 1518 3242 1521 3268
rect 1512 3203 1514 3207
rect 1518 3203 1521 3207
rect 1525 3203 1528 3207
rect 1398 3122 1401 3128
rect 1406 3092 1409 3128
rect 1430 3092 1433 3148
rect 1442 3138 1446 3141
rect 1462 3102 1465 3128
rect 1462 3092 1465 3098
rect 1494 3092 1497 3148
rect 1510 3142 1513 3178
rect 1518 3142 1521 3148
rect 1438 3078 1446 3081
rect 1506 3078 1510 3081
rect 1118 3032 1121 3038
rect 974 2992 977 3018
rect 850 2948 854 2951
rect 870 2942 873 2958
rect 918 2952 921 2978
rect 830 2938 838 2941
rect 834 2928 838 2931
rect 690 2878 694 2881
rect 718 2878 742 2881
rect 786 2878 790 2881
rect 654 2872 657 2878
rect 670 2872 673 2878
rect 718 2872 721 2878
rect 730 2868 734 2871
rect 638 2862 641 2868
rect 766 2862 769 2868
rect 774 2862 777 2868
rect 790 2862 793 2878
rect 806 2872 809 2928
rect 878 2921 881 2948
rect 926 2932 929 2938
rect 890 2928 894 2931
rect 914 2928 918 2931
rect 878 2918 889 2921
rect 854 2892 857 2918
rect 830 2882 833 2888
rect 818 2878 822 2881
rect 710 2852 713 2858
rect 718 2852 721 2858
rect 670 2842 673 2848
rect 638 2802 641 2818
rect 654 2792 657 2808
rect 638 2742 641 2768
rect 666 2748 670 2751
rect 678 2742 681 2798
rect 686 2792 689 2848
rect 718 2752 721 2828
rect 726 2812 729 2828
rect 694 2732 697 2738
rect 702 2732 705 2748
rect 726 2742 729 2808
rect 758 2742 761 2748
rect 766 2742 769 2748
rect 658 2728 662 2731
rect 714 2728 718 2731
rect 738 2728 742 2731
rect 614 2692 617 2698
rect 630 2671 633 2718
rect 686 2702 689 2718
rect 662 2698 670 2701
rect 638 2672 641 2678
rect 654 2672 657 2698
rect 662 2692 665 2698
rect 630 2668 638 2671
rect 550 2642 553 2648
rect 582 2642 585 2658
rect 606 2652 609 2668
rect 626 2658 630 2661
rect 650 2658 654 2661
rect 598 2642 601 2648
rect 602 2638 609 2641
rect 594 2628 601 2631
rect 482 2538 486 2541
rect 558 2532 561 2598
rect 566 2572 569 2618
rect 598 2592 601 2628
rect 582 2562 585 2568
rect 566 2552 569 2558
rect 590 2552 593 2558
rect 606 2541 609 2638
rect 614 2592 617 2648
rect 670 2631 673 2678
rect 678 2642 681 2678
rect 694 2672 697 2678
rect 702 2662 705 2708
rect 726 2682 729 2708
rect 774 2682 777 2758
rect 782 2752 785 2818
rect 798 2802 801 2818
rect 806 2802 809 2868
rect 814 2862 817 2868
rect 838 2852 841 2888
rect 862 2862 865 2868
rect 850 2858 854 2861
rect 870 2822 873 2868
rect 878 2862 881 2878
rect 782 2742 785 2748
rect 790 2742 793 2768
rect 822 2752 825 2768
rect 814 2742 817 2748
rect 802 2738 806 2741
rect 830 2741 833 2788
rect 846 2762 849 2818
rect 822 2738 833 2741
rect 854 2761 857 2818
rect 886 2782 889 2918
rect 894 2862 897 2918
rect 902 2882 905 2928
rect 934 2882 937 2988
rect 942 2952 945 2978
rect 950 2942 953 2958
rect 990 2942 993 2948
rect 1014 2942 1017 2948
rect 1022 2942 1025 2958
rect 1038 2942 1041 3018
rect 1062 2952 1065 2958
rect 1046 2942 1049 2948
rect 1078 2942 1081 2948
rect 1062 2938 1070 2941
rect 966 2932 969 2938
rect 974 2932 977 2938
rect 1050 2928 1054 2931
rect 982 2892 985 2918
rect 992 2903 994 2907
rect 998 2903 1001 2907
rect 1005 2903 1008 2907
rect 1022 2892 1025 2908
rect 1030 2902 1033 2918
rect 1046 2892 1049 2918
rect 926 2878 934 2881
rect 906 2868 910 2871
rect 926 2862 929 2878
rect 938 2868 942 2871
rect 910 2842 913 2848
rect 926 2832 929 2838
rect 854 2758 862 2761
rect 838 2742 841 2758
rect 846 2742 849 2758
rect 810 2728 817 2731
rect 754 2678 758 2681
rect 790 2678 798 2681
rect 734 2662 737 2668
rect 758 2662 761 2668
rect 770 2658 774 2661
rect 702 2642 705 2648
rect 686 2632 689 2638
rect 718 2632 721 2648
rect 670 2628 681 2631
rect 646 2582 649 2588
rect 622 2552 625 2558
rect 598 2538 609 2541
rect 614 2542 617 2548
rect 406 2522 409 2528
rect 502 2522 505 2528
rect 442 2518 446 2521
rect 458 2518 462 2521
rect 374 2422 377 2468
rect 406 2462 409 2488
rect 466 2478 470 2481
rect 446 2472 449 2478
rect 494 2472 497 2478
rect 522 2468 526 2471
rect 438 2462 441 2468
rect 518 2462 521 2468
rect 286 2362 289 2368
rect 278 2358 286 2361
rect 278 2332 281 2358
rect 302 2332 305 2338
rect 278 2262 281 2278
rect 246 2142 249 2148
rect 254 2132 257 2138
rect 262 2132 265 2218
rect 270 2162 273 2198
rect 278 2162 281 2168
rect 166 1952 169 1968
rect 174 1962 177 2018
rect 190 1971 193 2048
rect 182 1968 193 1971
rect 214 2002 217 2058
rect 238 2021 241 2078
rect 262 2072 265 2118
rect 278 2082 281 2118
rect 286 2082 289 2268
rect 294 2172 297 2318
rect 302 2262 305 2328
rect 310 2272 313 2398
rect 318 2372 321 2378
rect 342 2372 345 2378
rect 358 2372 361 2418
rect 374 2372 377 2418
rect 398 2392 401 2418
rect 406 2372 409 2458
rect 414 2432 417 2458
rect 474 2448 478 2451
rect 422 2442 425 2448
rect 502 2442 505 2448
rect 438 2382 441 2418
rect 334 2332 337 2338
rect 342 2331 345 2348
rect 342 2328 350 2331
rect 330 2278 334 2281
rect 302 2252 305 2258
rect 302 2152 305 2248
rect 310 2172 313 2268
rect 342 2252 345 2268
rect 334 2242 337 2248
rect 342 2162 345 2178
rect 310 2142 313 2158
rect 334 2152 337 2158
rect 302 2082 305 2088
rect 310 2072 313 2078
rect 318 2072 321 2148
rect 326 2112 329 2138
rect 334 2128 342 2131
rect 274 2068 278 2071
rect 246 2052 249 2068
rect 318 2062 321 2068
rect 262 2042 265 2058
rect 334 2052 337 2128
rect 350 2122 353 2308
rect 358 2292 361 2358
rect 366 2332 369 2358
rect 406 2342 409 2348
rect 394 2338 398 2341
rect 418 2338 422 2341
rect 442 2338 446 2341
rect 382 2332 385 2338
rect 414 2332 417 2338
rect 362 2268 366 2271
rect 374 2251 377 2318
rect 382 2262 385 2328
rect 402 2318 406 2321
rect 390 2272 393 2278
rect 414 2272 417 2328
rect 394 2268 401 2271
rect 370 2248 377 2251
rect 398 2252 401 2268
rect 430 2252 433 2328
rect 438 2312 441 2318
rect 442 2268 446 2271
rect 454 2261 457 2418
rect 462 2402 465 2438
rect 486 2422 489 2428
rect 480 2403 482 2407
rect 486 2403 489 2407
rect 493 2403 496 2407
rect 462 2362 465 2388
rect 502 2362 505 2418
rect 462 2272 465 2358
rect 442 2258 457 2261
rect 470 2261 473 2338
rect 482 2328 486 2331
rect 466 2258 473 2261
rect 494 2302 497 2308
rect 494 2262 497 2298
rect 502 2272 505 2358
rect 510 2352 513 2458
rect 542 2452 545 2508
rect 566 2492 569 2538
rect 574 2512 577 2518
rect 582 2471 585 2508
rect 574 2468 585 2471
rect 598 2482 601 2538
rect 670 2532 673 2538
rect 606 2522 609 2528
rect 630 2502 633 2528
rect 678 2522 681 2628
rect 686 2592 689 2608
rect 750 2602 753 2658
rect 770 2648 777 2651
rect 774 2642 777 2648
rect 750 2592 753 2598
rect 702 2532 705 2558
rect 718 2552 721 2568
rect 726 2562 729 2568
rect 734 2552 737 2558
rect 710 2542 713 2548
rect 758 2542 761 2628
rect 782 2612 785 2658
rect 790 2632 793 2678
rect 802 2658 806 2661
rect 806 2642 809 2648
rect 814 2622 817 2728
rect 822 2651 825 2738
rect 834 2728 838 2731
rect 854 2731 857 2748
rect 870 2742 873 2748
rect 886 2742 889 2748
rect 894 2742 897 2818
rect 910 2752 913 2778
rect 934 2772 937 2858
rect 950 2851 953 2888
rect 1034 2878 1038 2881
rect 982 2872 985 2878
rect 1054 2872 1057 2878
rect 1062 2872 1065 2938
rect 1074 2928 1078 2931
rect 1070 2882 1073 2888
rect 1018 2868 1025 2871
rect 966 2862 969 2868
rect 946 2848 953 2851
rect 950 2832 953 2848
rect 998 2792 1001 2858
rect 990 2772 993 2788
rect 946 2768 950 2771
rect 946 2758 950 2761
rect 1010 2758 1014 2761
rect 994 2748 998 2751
rect 846 2728 857 2731
rect 930 2738 934 2741
rect 862 2731 865 2738
rect 862 2728 886 2731
rect 838 2692 841 2698
rect 830 2662 833 2678
rect 846 2672 849 2728
rect 894 2701 897 2718
rect 894 2698 902 2701
rect 878 2691 881 2698
rect 878 2688 897 2691
rect 894 2681 897 2688
rect 870 2678 889 2681
rect 894 2678 905 2681
rect 822 2648 841 2651
rect 766 2552 769 2608
rect 794 2588 798 2591
rect 822 2572 825 2638
rect 838 2621 841 2648
rect 846 2632 849 2668
rect 854 2642 857 2658
rect 870 2652 873 2678
rect 886 2671 889 2678
rect 886 2668 894 2671
rect 870 2632 873 2648
rect 878 2642 881 2668
rect 902 2662 905 2678
rect 910 2662 913 2738
rect 918 2732 921 2738
rect 926 2702 929 2718
rect 930 2688 934 2691
rect 942 2672 945 2748
rect 950 2672 953 2708
rect 938 2658 942 2661
rect 918 2642 921 2648
rect 926 2642 929 2648
rect 838 2618 854 2621
rect 878 2612 881 2638
rect 886 2632 889 2638
rect 906 2628 910 2631
rect 830 2592 833 2598
rect 878 2592 881 2598
rect 958 2592 961 2748
rect 978 2738 982 2741
rect 992 2703 994 2707
rect 998 2703 1001 2707
rect 1005 2703 1008 2707
rect 1022 2692 1025 2868
rect 1030 2852 1033 2868
rect 1030 2732 1033 2828
rect 1062 2751 1065 2868
rect 1070 2862 1073 2868
rect 1086 2862 1089 2998
rect 1094 2952 1097 2958
rect 1102 2942 1105 2958
rect 1102 2932 1105 2938
rect 1110 2892 1113 3018
rect 1118 2992 1121 3028
rect 1222 3022 1225 3038
rect 1138 2958 1142 2961
rect 1118 2952 1121 2958
rect 1158 2952 1161 2958
rect 1130 2938 1134 2941
rect 1150 2902 1153 2938
rect 1110 2881 1113 2888
rect 1106 2878 1113 2881
rect 1098 2868 1102 2871
rect 1110 2851 1113 2868
rect 1118 2862 1121 2898
rect 1158 2892 1161 2908
rect 1166 2892 1169 2938
rect 1174 2932 1177 2938
rect 1182 2932 1185 2968
rect 1190 2942 1193 2948
rect 1214 2942 1217 2958
rect 1222 2952 1225 2978
rect 1198 2892 1201 2938
rect 1222 2932 1225 2938
rect 1230 2932 1233 3008
rect 1238 2992 1241 3068
rect 1246 3052 1249 3058
rect 1270 3052 1273 3058
rect 1310 3052 1313 3058
rect 1246 2988 1254 2991
rect 1246 2952 1249 2988
rect 1278 2961 1281 3018
rect 1258 2958 1265 2961
rect 1278 2958 1286 2961
rect 1210 2928 1214 2931
rect 1222 2892 1225 2928
rect 1134 2862 1137 2888
rect 1230 2882 1233 2928
rect 1238 2882 1241 2918
rect 1142 2862 1145 2868
rect 1110 2848 1121 2851
rect 1078 2842 1081 2848
rect 1118 2822 1121 2848
rect 1098 2788 1102 2791
rect 1062 2748 1070 2751
rect 1054 2722 1057 2728
rect 1062 2722 1065 2738
rect 1046 2692 1049 2708
rect 982 2622 985 2678
rect 1014 2642 1017 2668
rect 1030 2612 1033 2678
rect 1070 2671 1073 2748
rect 1086 2712 1089 2768
rect 1094 2742 1097 2748
rect 1102 2732 1105 2758
rect 1110 2742 1113 2808
rect 1118 2792 1121 2818
rect 1134 2812 1137 2818
rect 1134 2792 1137 2798
rect 1130 2758 1137 2761
rect 1094 2672 1097 2688
rect 1102 2678 1110 2681
rect 1070 2668 1078 2671
rect 1038 2652 1041 2658
rect 1054 2632 1057 2668
rect 1062 2652 1065 2658
rect 782 2562 785 2568
rect 786 2548 790 2551
rect 806 2542 809 2558
rect 830 2552 833 2578
rect 902 2562 905 2578
rect 1070 2562 1073 2618
rect 1078 2572 1081 2608
rect 1086 2592 1089 2658
rect 1102 2622 1105 2678
rect 1110 2662 1113 2668
rect 1118 2652 1121 2718
rect 1126 2662 1129 2748
rect 1134 2672 1137 2758
rect 1142 2742 1145 2848
rect 1150 2802 1153 2878
rect 1206 2872 1209 2878
rect 1230 2872 1233 2878
rect 1246 2872 1249 2948
rect 1254 2942 1257 2948
rect 1262 2932 1265 2958
rect 1270 2938 1278 2941
rect 1270 2882 1273 2938
rect 1278 2882 1281 2888
rect 1258 2878 1262 2881
rect 1286 2872 1289 2958
rect 1294 2892 1297 3048
rect 1310 3032 1313 3038
rect 1302 2972 1305 3008
rect 1310 2961 1313 3018
rect 1302 2958 1313 2961
rect 1318 2962 1321 2968
rect 1302 2942 1305 2958
rect 1310 2942 1313 2948
rect 1326 2942 1329 3048
rect 1342 3002 1345 3068
rect 1374 3062 1377 3078
rect 1366 3052 1369 3058
rect 1178 2868 1182 2871
rect 1302 2862 1305 2938
rect 1326 2922 1329 2928
rect 1318 2872 1321 2918
rect 1334 2892 1337 2958
rect 1342 2932 1345 2998
rect 1350 2972 1353 2978
rect 1358 2962 1361 3018
rect 1366 2972 1369 3048
rect 1378 3028 1382 3031
rect 1390 3022 1393 3078
rect 1398 3052 1401 3078
rect 1414 3052 1417 3068
rect 1350 2932 1353 2948
rect 1358 2942 1361 2958
rect 1366 2931 1369 2968
rect 1414 2962 1417 3048
rect 1422 3022 1425 3058
rect 1430 3042 1433 3058
rect 1438 3032 1441 3078
rect 1450 3048 1454 3051
rect 1430 3002 1433 3018
rect 1470 3002 1473 3068
rect 1478 3052 1481 3058
rect 1486 3052 1489 3068
rect 1526 3062 1529 3088
rect 1478 2992 1481 3018
rect 1450 2978 1454 2981
rect 1478 2972 1481 2988
rect 1442 2958 1446 2961
rect 1358 2928 1369 2931
rect 1358 2892 1361 2928
rect 1374 2922 1377 2928
rect 1326 2862 1329 2868
rect 1174 2852 1177 2858
rect 1198 2852 1201 2858
rect 1230 2852 1233 2858
rect 1270 2852 1273 2858
rect 1310 2852 1313 2858
rect 1218 2848 1222 2851
rect 1350 2851 1353 2878
rect 1366 2862 1369 2918
rect 1398 2872 1401 2938
rect 1422 2922 1425 2948
rect 1430 2942 1433 2958
rect 1454 2942 1457 2958
rect 1406 2912 1409 2918
rect 1406 2882 1409 2908
rect 1414 2892 1417 2908
rect 1430 2872 1433 2938
rect 1458 2928 1462 2931
rect 1378 2868 1382 2871
rect 1378 2858 1382 2861
rect 1406 2852 1409 2868
rect 1346 2848 1353 2851
rect 1198 2792 1201 2838
rect 1214 2762 1217 2848
rect 1270 2842 1273 2848
rect 1290 2838 1294 2841
rect 1270 2802 1273 2818
rect 1298 2788 1302 2791
rect 1150 2752 1153 2758
rect 1198 2752 1201 2758
rect 1178 2748 1182 2751
rect 1230 2751 1233 2758
rect 1214 2742 1217 2748
rect 1162 2738 1169 2741
rect 1142 2702 1145 2738
rect 1166 2692 1169 2738
rect 1174 2732 1177 2738
rect 1186 2728 1190 2731
rect 1222 2682 1225 2698
rect 1230 2692 1233 2708
rect 1174 2672 1177 2678
rect 1162 2668 1166 2671
rect 1134 2662 1137 2668
rect 1150 2662 1153 2668
rect 1210 2658 1214 2661
rect 1182 2652 1185 2658
rect 1230 2652 1233 2688
rect 1238 2672 1241 2768
rect 1242 2658 1246 2661
rect 1254 2651 1257 2698
rect 1286 2692 1289 2788
rect 1310 2742 1313 2848
rect 1350 2812 1353 2848
rect 1394 2848 1398 2851
rect 1302 2732 1305 2738
rect 1318 2732 1321 2748
rect 1326 2732 1329 2758
rect 1350 2752 1353 2778
rect 1338 2738 1342 2741
rect 1338 2728 1342 2731
rect 1262 2670 1265 2688
rect 1270 2672 1273 2678
rect 1246 2648 1257 2651
rect 1138 2638 1142 2641
rect 842 2558 846 2561
rect 874 2558 878 2561
rect 1110 2552 1113 2558
rect 1118 2552 1121 2638
rect 1126 2552 1129 2618
rect 1182 2592 1185 2648
rect 1210 2628 1214 2631
rect 1142 2552 1145 2588
rect 1190 2562 1193 2618
rect 1170 2558 1174 2561
rect 938 2548 942 2551
rect 970 2548 974 2551
rect 1018 2548 1022 2551
rect 918 2542 921 2548
rect 754 2538 758 2541
rect 930 2538 934 2541
rect 690 2528 694 2531
rect 598 2472 601 2478
rect 566 2462 569 2468
rect 574 2462 577 2468
rect 570 2448 574 2451
rect 534 2442 537 2448
rect 558 2402 561 2418
rect 582 2402 585 2458
rect 510 2342 513 2348
rect 530 2338 534 2341
rect 522 2328 526 2331
rect 462 2252 465 2258
rect 358 2212 361 2248
rect 366 2162 369 2168
rect 390 2162 393 2238
rect 406 2162 409 2218
rect 386 2148 390 2151
rect 362 2138 366 2141
rect 410 2138 414 2141
rect 342 2082 345 2118
rect 342 2072 345 2078
rect 350 2042 353 2058
rect 266 2038 273 2041
rect 238 2018 246 2021
rect 134 1888 142 1891
rect 110 1752 113 1758
rect 78 1742 81 1748
rect 86 1742 89 1748
rect 58 1648 65 1651
rect 54 1562 57 1568
rect 46 1548 57 1551
rect 54 1542 57 1548
rect 34 1538 38 1541
rect 6 1362 9 1478
rect 22 1462 25 1538
rect 22 1342 25 1458
rect 46 1452 49 1518
rect 54 1472 57 1538
rect 70 1531 73 1618
rect 78 1562 81 1698
rect 94 1671 97 1748
rect 118 1742 121 1858
rect 134 1762 137 1888
rect 142 1882 145 1888
rect 150 1872 153 1948
rect 174 1942 177 1948
rect 182 1942 185 1968
rect 190 1952 193 1958
rect 206 1952 209 1958
rect 162 1928 166 1931
rect 214 1912 217 1998
rect 230 1942 233 1988
rect 238 1952 241 1968
rect 246 1962 249 2018
rect 262 2012 265 2018
rect 210 1878 214 1881
rect 222 1872 225 1918
rect 150 1842 153 1868
rect 170 1848 174 1851
rect 142 1762 145 1778
rect 158 1752 161 1758
rect 162 1738 166 1741
rect 110 1682 113 1718
rect 118 1711 121 1738
rect 150 1722 153 1738
rect 174 1732 177 1748
rect 130 1718 134 1721
rect 118 1708 129 1711
rect 126 1692 129 1708
rect 182 1672 185 1858
rect 190 1792 193 1858
rect 190 1762 193 1788
rect 206 1762 209 1868
rect 230 1862 233 1928
rect 250 1918 254 1921
rect 222 1832 225 1858
rect 246 1852 249 1858
rect 254 1792 257 1858
rect 254 1762 257 1768
rect 198 1742 201 1748
rect 222 1712 225 1748
rect 238 1742 241 1748
rect 262 1742 265 1978
rect 270 1952 273 2038
rect 278 1952 281 2018
rect 286 1962 289 1988
rect 294 1982 297 2018
rect 274 1938 278 1941
rect 302 1932 305 1988
rect 310 1952 313 1978
rect 270 1852 273 1868
rect 286 1762 289 1918
rect 294 1872 297 1918
rect 318 1902 321 2018
rect 338 1948 342 1951
rect 350 1942 353 1948
rect 314 1858 318 1861
rect 294 1842 297 1858
rect 294 1762 297 1838
rect 270 1752 273 1758
rect 294 1742 297 1758
rect 230 1732 233 1738
rect 242 1688 246 1691
rect 254 1682 257 1718
rect 90 1668 97 1671
rect 86 1562 89 1638
rect 94 1562 97 1668
rect 218 1668 222 1671
rect 110 1652 113 1658
rect 158 1652 161 1658
rect 102 1642 105 1648
rect 166 1632 169 1668
rect 210 1658 214 1661
rect 222 1652 225 1658
rect 186 1648 190 1651
rect 150 1612 153 1618
rect 102 1552 105 1558
rect 126 1552 129 1588
rect 150 1562 153 1568
rect 138 1558 142 1561
rect 154 1558 158 1561
rect 146 1548 150 1551
rect 118 1542 121 1548
rect 70 1528 81 1531
rect 54 1441 57 1468
rect 46 1438 57 1441
rect 30 1362 33 1418
rect 46 1352 49 1438
rect 62 1432 65 1438
rect 70 1372 73 1518
rect 78 1492 81 1528
rect 94 1482 97 1538
rect 126 1472 129 1548
rect 166 1542 169 1618
rect 190 1562 193 1568
rect 198 1552 201 1648
rect 230 1642 233 1658
rect 206 1632 209 1638
rect 218 1578 222 1581
rect 230 1552 233 1638
rect 238 1552 241 1678
rect 262 1672 265 1738
rect 258 1658 262 1661
rect 270 1652 273 1678
rect 210 1548 214 1551
rect 198 1542 201 1548
rect 154 1528 158 1531
rect 166 1522 169 1538
rect 174 1532 177 1538
rect 174 1472 177 1478
rect 98 1468 102 1471
rect 98 1458 102 1461
rect 78 1452 81 1458
rect 98 1448 102 1451
rect 114 1448 118 1451
rect 126 1442 129 1468
rect 54 1362 57 1368
rect 86 1352 89 1418
rect 102 1362 105 1368
rect 110 1352 113 1358
rect 46 1342 49 1348
rect 26 1338 30 1341
rect 14 1312 17 1318
rect 14 1282 17 1288
rect 14 1192 17 1258
rect 30 1252 33 1258
rect 38 1161 41 1318
rect 54 1261 57 1318
rect 62 1292 65 1308
rect 70 1292 73 1348
rect 134 1342 137 1458
rect 166 1452 169 1458
rect 182 1452 185 1518
rect 190 1462 193 1528
rect 206 1472 209 1478
rect 198 1462 201 1468
rect 194 1458 198 1461
rect 146 1448 150 1451
rect 166 1422 169 1438
rect 166 1362 169 1418
rect 182 1362 185 1368
rect 142 1342 145 1348
rect 166 1342 169 1348
rect 190 1342 193 1348
rect 90 1338 94 1341
rect 130 1338 134 1341
rect 50 1258 57 1261
rect 66 1258 70 1261
rect 70 1232 73 1258
rect 78 1212 81 1258
rect 86 1252 89 1258
rect 94 1172 97 1318
rect 110 1262 113 1328
rect 130 1278 134 1281
rect 34 1158 41 1161
rect 62 1162 65 1168
rect 102 1162 105 1218
rect 78 1158 86 1161
rect 90 1158 94 1161
rect 6 1132 9 1138
rect 6 1092 9 1118
rect 14 1062 17 1148
rect 30 1061 33 1148
rect 42 1138 46 1141
rect 54 1082 57 1138
rect 70 1132 73 1138
rect 78 1132 81 1158
rect 102 1142 105 1148
rect 110 1142 113 1258
rect 126 1162 129 1278
rect 134 1252 137 1258
rect 134 1192 137 1248
rect 142 1192 145 1218
rect 150 1161 153 1318
rect 166 1282 169 1288
rect 162 1268 166 1271
rect 166 1162 169 1168
rect 150 1158 158 1161
rect 174 1161 177 1318
rect 198 1282 201 1418
rect 214 1362 217 1548
rect 254 1531 257 1568
rect 270 1562 273 1608
rect 246 1528 257 1531
rect 262 1532 265 1558
rect 246 1462 249 1528
rect 254 1502 257 1518
rect 222 1442 225 1458
rect 254 1452 257 1458
rect 270 1451 273 1518
rect 278 1462 281 1738
rect 302 1731 305 1858
rect 310 1762 313 1818
rect 294 1728 305 1731
rect 286 1702 289 1718
rect 294 1672 297 1728
rect 318 1722 321 1728
rect 310 1682 313 1718
rect 302 1672 305 1678
rect 286 1572 289 1618
rect 294 1602 297 1658
rect 310 1622 313 1658
rect 318 1642 321 1718
rect 326 1682 329 1918
rect 334 1862 337 1898
rect 350 1872 353 1938
rect 334 1722 337 1728
rect 326 1652 329 1668
rect 342 1662 345 1868
rect 350 1842 353 1868
rect 358 1851 361 2058
rect 366 2052 369 2118
rect 382 2062 385 2098
rect 390 2062 393 2138
rect 406 2062 409 2128
rect 374 2002 377 2058
rect 374 1962 377 1988
rect 382 1952 385 1958
rect 398 1952 401 2018
rect 394 1938 398 1941
rect 406 1922 409 1938
rect 366 1872 369 1918
rect 382 1862 385 1898
rect 358 1848 366 1851
rect 358 1772 361 1818
rect 366 1761 369 1848
rect 374 1842 377 1858
rect 390 1792 393 1918
rect 414 1902 417 2118
rect 422 2082 425 2218
rect 430 2152 433 2168
rect 446 2152 449 2208
rect 446 2142 449 2148
rect 454 2112 457 2148
rect 462 2112 465 2248
rect 480 2203 482 2207
rect 486 2203 489 2207
rect 493 2203 496 2207
rect 478 2162 481 2168
rect 438 2072 441 2078
rect 422 1992 425 2008
rect 430 1992 433 2018
rect 422 1962 425 1988
rect 430 1962 433 1978
rect 438 1962 441 2068
rect 446 2042 449 2068
rect 454 2062 457 2098
rect 470 2092 473 2118
rect 446 1942 449 1948
rect 422 1881 425 1918
rect 454 1902 457 1918
rect 414 1878 425 1881
rect 382 1762 385 1768
rect 362 1758 369 1761
rect 350 1752 353 1758
rect 374 1742 377 1758
rect 398 1752 401 1838
rect 414 1762 417 1878
rect 422 1822 425 1868
rect 430 1862 433 1898
rect 462 1871 465 2028
rect 470 1922 473 2068
rect 478 2052 481 2118
rect 494 2062 497 2068
rect 502 2032 505 2218
rect 510 2152 513 2318
rect 518 2262 521 2268
rect 526 2252 529 2258
rect 534 2252 537 2318
rect 542 2292 545 2358
rect 550 2352 553 2358
rect 566 2322 569 2348
rect 582 2342 585 2378
rect 590 2352 593 2448
rect 590 2331 593 2348
rect 598 2342 601 2458
rect 606 2452 609 2478
rect 622 2462 625 2468
rect 630 2451 633 2498
rect 662 2472 665 2478
rect 674 2458 678 2461
rect 622 2448 633 2451
rect 686 2452 689 2458
rect 710 2452 713 2488
rect 742 2472 745 2528
rect 766 2482 769 2538
rect 774 2492 777 2518
rect 802 2498 809 2501
rect 778 2468 782 2471
rect 806 2462 809 2498
rect 830 2462 833 2528
rect 846 2512 849 2538
rect 894 2532 897 2538
rect 866 2528 870 2531
rect 870 2522 873 2528
rect 754 2458 758 2461
rect 826 2458 830 2461
rect 614 2372 617 2418
rect 614 2342 617 2358
rect 582 2328 593 2331
rect 614 2332 617 2338
rect 550 2302 553 2318
rect 570 2278 574 2281
rect 582 2272 585 2328
rect 606 2312 609 2318
rect 594 2278 598 2281
rect 614 2281 617 2308
rect 610 2278 617 2281
rect 550 2262 553 2268
rect 558 2222 561 2268
rect 574 2252 577 2268
rect 614 2262 617 2268
rect 622 2262 625 2448
rect 674 2418 678 2421
rect 638 2362 641 2368
rect 630 2302 633 2358
rect 646 2331 649 2418
rect 694 2392 697 2418
rect 710 2402 713 2448
rect 726 2392 729 2458
rect 766 2452 769 2458
rect 790 2452 793 2458
rect 750 2382 753 2418
rect 758 2372 761 2398
rect 702 2362 705 2368
rect 734 2362 737 2368
rect 666 2358 670 2361
rect 754 2358 758 2361
rect 674 2348 678 2351
rect 654 2342 657 2348
rect 686 2342 689 2348
rect 666 2338 670 2341
rect 646 2328 657 2331
rect 642 2318 646 2321
rect 646 2252 649 2258
rect 590 2242 593 2248
rect 550 2172 553 2218
rect 582 2202 585 2218
rect 546 2158 550 2161
rect 518 2112 521 2138
rect 518 2072 521 2088
rect 526 2062 529 2068
rect 526 2012 529 2018
rect 480 2003 482 2007
rect 486 2003 489 2007
rect 493 2003 496 2007
rect 478 1952 481 1978
rect 502 1962 505 1998
rect 478 1932 481 1938
rect 502 1912 505 1918
rect 510 1882 513 2008
rect 534 2002 537 2118
rect 542 2052 545 2118
rect 550 2062 553 2088
rect 558 2082 561 2148
rect 566 2142 569 2188
rect 630 2171 633 2218
rect 654 2202 657 2328
rect 666 2278 670 2281
rect 678 2272 681 2308
rect 686 2272 689 2338
rect 694 2312 697 2338
rect 706 2318 710 2321
rect 718 2321 721 2348
rect 726 2342 729 2358
rect 766 2342 769 2438
rect 774 2352 777 2368
rect 790 2362 793 2378
rect 786 2348 790 2351
rect 802 2348 806 2351
rect 814 2342 817 2448
rect 838 2442 841 2458
rect 854 2451 857 2518
rect 878 2481 881 2518
rect 870 2478 881 2481
rect 870 2472 873 2478
rect 878 2462 881 2468
rect 850 2448 857 2451
rect 822 2362 825 2418
rect 846 2362 849 2448
rect 858 2418 862 2421
rect 854 2362 857 2378
rect 870 2352 873 2458
rect 886 2452 889 2518
rect 894 2452 897 2528
rect 910 2472 913 2518
rect 902 2462 905 2468
rect 934 2462 937 2468
rect 922 2458 926 2461
rect 922 2448 926 2451
rect 886 2382 889 2418
rect 910 2372 913 2418
rect 942 2411 945 2548
rect 954 2538 958 2541
rect 1002 2538 1006 2541
rect 1042 2538 1046 2541
rect 1074 2538 1078 2541
rect 1090 2540 1094 2543
rect 1174 2542 1177 2548
rect 1130 2538 1134 2541
rect 1146 2538 1150 2541
rect 950 2452 953 2518
rect 958 2462 961 2528
rect 982 2492 985 2518
rect 1030 2512 1033 2518
rect 992 2503 994 2507
rect 998 2503 1001 2507
rect 1005 2503 1008 2507
rect 1038 2472 1041 2518
rect 1054 2492 1057 2538
rect 1106 2518 1110 2521
rect 1062 2502 1065 2518
rect 1118 2492 1121 2538
rect 1130 2528 1134 2531
rect 1174 2512 1177 2528
rect 1198 2522 1201 2558
rect 1214 2552 1217 2558
rect 1230 2542 1233 2628
rect 1238 2592 1241 2598
rect 1246 2542 1249 2648
rect 1278 2572 1281 2658
rect 1294 2592 1297 2728
rect 1350 2712 1353 2748
rect 1358 2742 1361 2798
rect 1374 2742 1377 2838
rect 1382 2752 1385 2848
rect 1390 2792 1393 2808
rect 1334 2692 1337 2708
rect 1290 2588 1294 2591
rect 1302 2572 1305 2658
rect 1318 2652 1321 2668
rect 1310 2602 1313 2618
rect 1318 2612 1321 2648
rect 1310 2582 1313 2598
rect 1334 2552 1337 2588
rect 1350 2582 1353 2658
rect 1358 2652 1361 2728
rect 1366 2662 1369 2718
rect 1382 2682 1385 2748
rect 1398 2742 1401 2758
rect 1406 2752 1409 2838
rect 1398 2692 1401 2728
rect 1406 2692 1409 2748
rect 1422 2742 1425 2868
rect 1438 2861 1441 2898
rect 1454 2882 1457 2898
rect 1434 2858 1441 2861
rect 1438 2842 1441 2858
rect 1462 2862 1465 2878
rect 1470 2872 1473 2968
rect 1494 2962 1497 2998
rect 1502 2962 1505 3008
rect 1512 3003 1514 3007
rect 1518 3003 1521 3007
rect 1525 3003 1528 3007
rect 1534 2962 1537 3328
rect 1550 3302 1553 3328
rect 1574 3272 1577 3328
rect 1598 3302 1601 3328
rect 1646 3302 1649 3328
rect 1670 3302 1673 3328
rect 1634 3288 1638 3291
rect 1566 3262 1569 3268
rect 1590 3262 1593 3278
rect 1654 3272 1657 3278
rect 1642 3268 1646 3271
rect 1670 3262 1673 3288
rect 1542 3102 1545 3238
rect 1566 3182 1569 3258
rect 1638 3252 1641 3258
rect 1574 3192 1577 3238
rect 1598 3172 1601 3218
rect 1678 3202 1681 3328
rect 1702 3282 1705 3328
rect 1726 3302 1729 3328
rect 1686 3252 1689 3278
rect 1702 3262 1705 3268
rect 1730 3258 1734 3261
rect 1598 3132 1601 3168
rect 1666 3148 1670 3151
rect 1542 3082 1545 3098
rect 1578 3088 1582 3091
rect 1590 3082 1593 3118
rect 1574 3078 1582 3081
rect 1542 3041 1545 3078
rect 1554 3048 1558 3051
rect 1566 3042 1569 3078
rect 1542 3038 1553 3041
rect 1550 3022 1553 3038
rect 1566 3002 1569 3038
rect 1522 2958 1526 2961
rect 1494 2932 1497 2958
rect 1534 2942 1537 2958
rect 1558 2952 1561 2988
rect 1574 2942 1577 3078
rect 1582 3052 1585 3068
rect 1582 2992 1585 3018
rect 1506 2918 1510 2921
rect 1490 2878 1497 2881
rect 1494 2872 1497 2878
rect 1482 2868 1486 2871
rect 1482 2858 1489 2861
rect 1498 2858 1502 2861
rect 1430 2762 1433 2838
rect 1462 2762 1465 2858
rect 1486 2792 1489 2858
rect 1526 2852 1529 2858
rect 1512 2803 1514 2807
rect 1518 2803 1521 2807
rect 1525 2803 1528 2807
rect 1430 2752 1433 2758
rect 1414 2712 1417 2718
rect 1422 2672 1425 2728
rect 1414 2652 1417 2658
rect 1354 2558 1358 2561
rect 1314 2548 1318 2551
rect 1366 2542 1369 2548
rect 1222 2532 1225 2538
rect 1002 2468 1006 2471
rect 1062 2462 1065 2478
rect 1126 2471 1129 2498
rect 1122 2468 1129 2471
rect 1154 2468 1158 2471
rect 1166 2462 1169 2488
rect 1002 2458 1006 2461
rect 1138 2458 1142 2461
rect 974 2442 977 2448
rect 966 2422 969 2438
rect 934 2408 945 2411
rect 918 2382 921 2388
rect 878 2358 886 2361
rect 822 2342 825 2348
rect 830 2342 833 2348
rect 786 2338 790 2341
rect 734 2322 737 2338
rect 854 2322 857 2328
rect 718 2318 726 2321
rect 762 2318 766 2321
rect 806 2282 809 2318
rect 794 2278 798 2281
rect 758 2272 761 2278
rect 766 2272 769 2278
rect 686 2262 689 2268
rect 710 2262 713 2268
rect 686 2252 689 2258
rect 750 2252 753 2258
rect 666 2238 670 2241
rect 690 2238 694 2241
rect 726 2212 729 2238
rect 758 2222 761 2268
rect 782 2232 785 2268
rect 822 2262 825 2288
rect 846 2282 849 2318
rect 862 2272 865 2348
rect 870 2322 873 2348
rect 878 2292 881 2358
rect 902 2352 905 2358
rect 890 2348 894 2351
rect 910 2342 913 2348
rect 934 2342 937 2408
rect 950 2362 953 2418
rect 942 2352 945 2358
rect 966 2342 969 2418
rect 982 2402 985 2458
rect 990 2412 993 2458
rect 1054 2452 1057 2458
rect 998 2362 1001 2438
rect 1002 2348 1006 2351
rect 974 2342 977 2348
rect 1014 2342 1017 2408
rect 1030 2362 1033 2398
rect 1038 2342 1041 2438
rect 1046 2402 1049 2418
rect 854 2262 857 2268
rect 846 2251 849 2258
rect 878 2252 881 2268
rect 846 2248 878 2251
rect 630 2168 638 2171
rect 678 2162 681 2168
rect 718 2162 721 2198
rect 590 2152 593 2158
rect 598 2152 601 2158
rect 622 2142 625 2148
rect 566 2132 569 2138
rect 602 2118 606 2121
rect 566 2052 569 2118
rect 574 2112 577 2118
rect 590 2072 593 2098
rect 606 2062 609 2068
rect 614 2062 617 2138
rect 622 2102 625 2138
rect 630 2132 633 2148
rect 630 2062 633 2098
rect 638 2082 641 2138
rect 646 2122 649 2158
rect 726 2152 729 2198
rect 750 2152 753 2218
rect 774 2162 777 2218
rect 798 2202 801 2218
rect 822 2162 825 2168
rect 838 2152 841 2218
rect 886 2202 889 2268
rect 894 2202 897 2338
rect 926 2331 929 2338
rect 926 2328 937 2331
rect 918 2281 921 2318
rect 910 2278 921 2281
rect 910 2272 913 2278
rect 918 2262 921 2268
rect 926 2262 929 2298
rect 934 2292 937 2328
rect 958 2312 961 2318
rect 1014 2312 1017 2338
rect 1046 2332 1049 2348
rect 992 2303 994 2307
rect 998 2303 1001 2307
rect 1005 2303 1008 2307
rect 950 2262 953 2278
rect 998 2262 1001 2288
rect 906 2258 910 2261
rect 974 2232 977 2258
rect 1006 2242 1009 2258
rect 854 2162 857 2168
rect 894 2162 897 2168
rect 690 2138 694 2141
rect 654 2132 657 2138
rect 702 2132 705 2138
rect 726 2132 729 2138
rect 758 2132 761 2138
rect 682 2118 686 2121
rect 642 2068 646 2071
rect 662 2061 665 2118
rect 674 2068 678 2071
rect 662 2058 673 2061
rect 550 1982 553 2018
rect 534 1962 537 1978
rect 526 1952 529 1958
rect 550 1952 553 1978
rect 558 1942 561 1968
rect 566 1962 569 1988
rect 562 1938 566 1941
rect 526 1932 529 1938
rect 526 1882 529 1908
rect 482 1878 486 1881
rect 454 1868 465 1871
rect 534 1872 537 1928
rect 454 1862 457 1868
rect 438 1772 441 1818
rect 454 1772 457 1858
rect 462 1852 465 1858
rect 534 1852 537 1858
rect 518 1832 521 1838
rect 470 1802 473 1818
rect 480 1803 482 1807
rect 486 1803 489 1807
rect 493 1803 496 1807
rect 426 1748 430 1751
rect 370 1738 374 1741
rect 426 1738 430 1741
rect 406 1732 409 1738
rect 438 1722 441 1738
rect 358 1672 361 1718
rect 382 1712 385 1718
rect 366 1662 369 1668
rect 390 1662 393 1678
rect 438 1662 441 1668
rect 418 1658 422 1661
rect 334 1652 337 1658
rect 306 1568 310 1571
rect 318 1562 321 1598
rect 334 1552 337 1598
rect 286 1532 289 1538
rect 294 1532 297 1538
rect 294 1481 297 1528
rect 286 1478 297 1481
rect 286 1472 289 1478
rect 302 1472 305 1548
rect 318 1542 321 1548
rect 298 1468 302 1471
rect 282 1458 286 1461
rect 266 1448 273 1451
rect 234 1438 238 1441
rect 230 1362 233 1388
rect 238 1362 241 1368
rect 254 1342 257 1348
rect 262 1342 265 1408
rect 186 1268 190 1271
rect 198 1262 201 1268
rect 186 1258 190 1261
rect 186 1248 190 1251
rect 198 1242 201 1248
rect 206 1172 209 1318
rect 214 1272 217 1338
rect 246 1332 249 1338
rect 266 1328 270 1331
rect 214 1262 217 1268
rect 222 1252 225 1258
rect 230 1252 233 1318
rect 254 1292 257 1318
rect 278 1282 281 1418
rect 294 1352 297 1468
rect 310 1452 313 1508
rect 318 1452 321 1538
rect 342 1522 345 1658
rect 354 1628 358 1631
rect 358 1552 361 1568
rect 362 1548 369 1551
rect 350 1512 353 1518
rect 326 1482 329 1508
rect 338 1478 342 1481
rect 330 1458 334 1461
rect 302 1381 305 1418
rect 310 1392 313 1448
rect 350 1432 353 1478
rect 358 1452 361 1458
rect 302 1378 313 1381
rect 250 1278 254 1281
rect 302 1272 305 1368
rect 310 1362 313 1378
rect 318 1372 321 1418
rect 342 1362 345 1378
rect 366 1362 369 1548
rect 374 1542 377 1658
rect 382 1602 385 1658
rect 430 1652 433 1658
rect 446 1622 449 1748
rect 454 1742 457 1748
rect 478 1702 481 1748
rect 490 1738 494 1741
rect 502 1732 505 1818
rect 526 1762 529 1828
rect 542 1821 545 1938
rect 550 1832 553 1858
rect 558 1852 561 1878
rect 566 1852 569 1918
rect 574 1912 577 2058
rect 590 2031 593 2058
rect 598 2042 601 2058
rect 582 2028 593 2031
rect 582 1962 585 2028
rect 590 1962 593 1988
rect 614 1962 617 2008
rect 622 1992 625 2018
rect 646 1962 649 2058
rect 654 2042 657 2058
rect 662 2042 665 2048
rect 654 2012 657 2018
rect 658 1988 662 1991
rect 670 1962 673 2058
rect 686 2052 689 2078
rect 710 2072 713 2128
rect 718 2071 721 2118
rect 750 2112 753 2118
rect 758 2092 761 2108
rect 718 2068 729 2071
rect 686 2042 689 2048
rect 694 2032 697 2068
rect 710 2062 713 2068
rect 650 1948 654 1951
rect 662 1951 665 1958
rect 662 1948 670 1951
rect 582 1942 585 1948
rect 606 1942 609 1948
rect 630 1942 633 1948
rect 638 1942 641 1948
rect 694 1942 697 1978
rect 710 1952 713 2058
rect 718 2042 721 2058
rect 726 1962 729 2068
rect 738 2058 742 2061
rect 750 2052 753 2078
rect 758 2072 761 2088
rect 758 2032 761 2068
rect 766 2062 769 2088
rect 774 2052 777 2148
rect 798 2142 801 2148
rect 918 2142 921 2188
rect 942 2172 945 2218
rect 958 2162 961 2198
rect 982 2162 985 2168
rect 950 2152 953 2158
rect 826 2138 830 2141
rect 882 2138 886 2141
rect 930 2138 934 2141
rect 978 2138 982 2141
rect 806 2132 809 2138
rect 782 2052 785 2118
rect 790 2082 793 2088
rect 734 1992 737 2018
rect 734 1962 737 1978
rect 590 1882 593 1918
rect 610 1878 614 1881
rect 582 1862 585 1868
rect 590 1852 593 1868
rect 614 1862 617 1868
rect 542 1818 553 1821
rect 526 1752 529 1758
rect 534 1742 537 1748
rect 542 1742 545 1768
rect 510 1732 513 1738
rect 502 1671 505 1728
rect 498 1668 505 1671
rect 506 1658 510 1661
rect 454 1652 457 1658
rect 494 1651 497 1658
rect 518 1652 521 1718
rect 534 1702 537 1718
rect 534 1672 537 1698
rect 550 1681 553 1818
rect 566 1752 569 1788
rect 558 1722 561 1728
rect 582 1712 585 1818
rect 590 1792 593 1828
rect 598 1802 601 1818
rect 606 1752 609 1818
rect 622 1782 625 1938
rect 646 1932 649 1938
rect 630 1852 633 1908
rect 630 1771 633 1848
rect 622 1768 633 1771
rect 622 1762 625 1768
rect 638 1761 641 1918
rect 646 1862 649 1928
rect 662 1872 665 1938
rect 742 1932 745 2028
rect 766 1992 769 2018
rect 770 1968 774 1971
rect 782 1962 785 1968
rect 790 1952 793 1988
rect 798 1972 801 2098
rect 806 2062 809 2128
rect 806 1992 809 2058
rect 822 2051 825 2118
rect 838 2102 841 2118
rect 838 2082 841 2088
rect 854 2082 857 2118
rect 862 2062 865 2138
rect 870 2112 873 2138
rect 918 2122 921 2138
rect 990 2121 993 2218
rect 1014 2172 1017 2258
rect 1030 2252 1033 2318
rect 1054 2302 1057 2338
rect 1046 2262 1049 2278
rect 1054 2272 1057 2278
rect 1062 2272 1065 2458
rect 1070 2362 1073 2408
rect 1078 2262 1081 2458
rect 1118 2452 1121 2458
rect 1090 2448 1094 2451
rect 1094 2362 1097 2438
rect 1110 2372 1113 2418
rect 1126 2402 1129 2448
rect 1142 2432 1145 2438
rect 1090 2338 1094 2341
rect 1102 2282 1105 2338
rect 1098 2268 1105 2271
rect 1082 2258 1086 2261
rect 1034 2248 1062 2251
rect 1070 2172 1073 2258
rect 1054 2162 1057 2168
rect 1078 2162 1081 2198
rect 1094 2172 1097 2258
rect 1102 2212 1105 2268
rect 1110 2152 1113 2348
rect 1118 2342 1121 2368
rect 1142 2362 1145 2368
rect 1150 2352 1153 2378
rect 1158 2372 1161 2458
rect 1166 2412 1169 2458
rect 1182 2442 1185 2518
rect 1206 2472 1209 2478
rect 1182 2412 1185 2418
rect 1190 2372 1193 2458
rect 1158 2352 1161 2368
rect 1190 2352 1193 2368
rect 1198 2342 1201 2458
rect 1206 2442 1209 2468
rect 1230 2462 1233 2538
rect 1238 2472 1241 2518
rect 1246 2492 1249 2538
rect 1254 2502 1257 2518
rect 1254 2472 1257 2478
rect 1262 2462 1265 2538
rect 1318 2532 1321 2538
rect 1242 2458 1246 2461
rect 1226 2448 1230 2451
rect 1270 2451 1273 2518
rect 1286 2472 1289 2508
rect 1326 2502 1329 2518
rect 1322 2488 1326 2491
rect 1294 2472 1297 2478
rect 1302 2462 1305 2468
rect 1358 2462 1361 2508
rect 1374 2502 1377 2638
rect 1382 2471 1385 2618
rect 1394 2568 1398 2571
rect 1406 2542 1409 2578
rect 1422 2572 1425 2658
rect 1430 2592 1433 2718
rect 1446 2712 1449 2748
rect 1454 2742 1457 2748
rect 1454 2672 1457 2738
rect 1462 2732 1465 2738
rect 1470 2712 1473 2748
rect 1486 2728 1494 2731
rect 1470 2672 1473 2688
rect 1486 2662 1489 2728
rect 1502 2722 1505 2728
rect 1510 2672 1513 2738
rect 1526 2731 1529 2788
rect 1534 2772 1537 2938
rect 1550 2922 1553 2938
rect 1566 2912 1569 2938
rect 1598 2932 1601 2958
rect 1562 2888 1566 2891
rect 1546 2878 1550 2881
rect 1570 2868 1574 2871
rect 1542 2772 1545 2818
rect 1574 2792 1577 2858
rect 1574 2772 1577 2778
rect 1538 2758 1542 2761
rect 1570 2748 1577 2751
rect 1526 2728 1534 2731
rect 1534 2692 1537 2728
rect 1498 2658 1502 2661
rect 1454 2652 1457 2658
rect 1454 2602 1457 2648
rect 1526 2642 1529 2678
rect 1534 2661 1537 2688
rect 1542 2672 1545 2748
rect 1566 2732 1569 2738
rect 1534 2658 1542 2661
rect 1550 2661 1553 2728
rect 1566 2672 1569 2728
rect 1574 2722 1577 2748
rect 1582 2742 1585 2888
rect 1598 2878 1601 2918
rect 1606 2912 1609 3138
rect 1638 3092 1641 3118
rect 1646 3092 1649 3108
rect 1654 3102 1657 3138
rect 1662 3122 1665 3128
rect 1670 3092 1673 3138
rect 1678 3132 1681 3188
rect 1686 3172 1689 3248
rect 1742 3182 1745 3328
rect 1790 3262 1793 3268
rect 1806 3252 1809 3278
rect 1818 3258 1822 3261
rect 1766 3232 1769 3238
rect 1778 3168 1782 3171
rect 1822 3162 1825 3168
rect 1730 3158 1734 3161
rect 1686 3152 1689 3158
rect 1698 3148 1702 3151
rect 1722 3148 1726 3151
rect 1738 3148 1742 3151
rect 1762 3148 1766 3151
rect 1718 3142 1721 3148
rect 1782 3142 1785 3148
rect 1738 3138 1742 3141
rect 1694 3132 1697 3138
rect 1806 3132 1809 3140
rect 1678 3122 1681 3128
rect 1618 3078 1622 3081
rect 1614 3072 1617 3078
rect 1662 3072 1665 3088
rect 1710 3082 1713 3088
rect 1678 3072 1681 3078
rect 1626 3068 1630 3071
rect 1630 3052 1633 3058
rect 1654 3052 1657 3058
rect 1646 3042 1649 3048
rect 1618 3038 1622 3041
rect 1614 2912 1617 2948
rect 1622 2932 1625 2938
rect 1630 2932 1633 2938
rect 1686 2932 1689 2958
rect 1694 2952 1697 3068
rect 1702 3062 1705 3068
rect 1702 2952 1705 3018
rect 1658 2918 1662 2921
rect 1630 2872 1633 2878
rect 1646 2872 1649 2908
rect 1694 2881 1697 2918
rect 1690 2878 1697 2881
rect 1710 2882 1713 3018
rect 1726 3012 1729 3058
rect 1726 2952 1729 2968
rect 1734 2951 1737 3038
rect 1742 2972 1745 3128
rect 1758 3122 1761 3128
rect 1758 3072 1761 3118
rect 1814 3112 1817 3138
rect 1766 2952 1769 3098
rect 1806 3072 1809 3108
rect 1814 3082 1817 3088
rect 1822 3082 1825 3148
rect 1830 3102 1833 3268
rect 1846 3262 1849 3268
rect 1838 3192 1841 3258
rect 1854 3222 1857 3258
rect 1846 3152 1849 3158
rect 1838 3112 1841 3148
rect 1846 3132 1849 3138
rect 1854 3132 1857 3168
rect 1826 3068 1830 3071
rect 1790 3062 1793 3068
rect 1774 2992 1777 3018
rect 1798 2992 1801 3058
rect 1846 3052 1849 3068
rect 1846 3042 1849 3048
rect 1862 3042 1865 3328
rect 1886 3328 1890 3332
rect 1950 3328 1954 3332
rect 1974 3328 1978 3332
rect 1990 3328 1994 3332
rect 2046 3331 2050 3332
rect 2094 3331 2098 3332
rect 2166 3331 2170 3332
rect 2046 3328 2057 3331
rect 2094 3328 2105 3331
rect 2166 3328 2177 3331
rect 1874 3248 1878 3251
rect 1870 3152 1873 3178
rect 1862 3022 1865 3028
rect 1774 2952 1777 2978
rect 1734 2948 1742 2951
rect 1718 2912 1721 2918
rect 1718 2872 1721 2908
rect 1726 2882 1729 2948
rect 1734 2872 1737 2938
rect 1766 2932 1769 2938
rect 1742 2922 1745 2928
rect 1746 2878 1750 2881
rect 1766 2872 1769 2878
rect 1774 2872 1777 2948
rect 1782 2942 1785 2958
rect 1822 2942 1825 2998
rect 1830 2952 1833 2998
rect 1838 2992 1841 3018
rect 1870 2982 1873 3128
rect 1878 3092 1881 3118
rect 1886 3082 1889 3328
rect 1950 3302 1953 3328
rect 1918 3272 1921 3278
rect 1894 3252 1897 3258
rect 1902 3252 1905 3268
rect 1902 3172 1905 3248
rect 1934 3232 1937 3268
rect 1954 3259 1958 3262
rect 1934 3162 1937 3228
rect 1974 3202 1977 3328
rect 1990 3302 1993 3328
rect 2024 3303 2026 3307
rect 2030 3303 2033 3307
rect 2037 3303 2040 3307
rect 2054 3292 2057 3328
rect 2102 3292 2105 3328
rect 2174 3292 2177 3328
rect 2230 3328 2234 3332
rect 2246 3328 2250 3332
rect 2262 3328 2266 3332
rect 2278 3331 2282 3332
rect 2270 3328 2282 3331
rect 2294 3328 2298 3332
rect 2310 3331 2314 3332
rect 2302 3328 2314 3331
rect 2326 3328 2330 3332
rect 2342 3331 2346 3332
rect 2414 3331 2418 3332
rect 2438 3331 2442 3332
rect 2342 3328 2353 3331
rect 2230 3302 2233 3328
rect 2246 3302 2249 3328
rect 2262 3302 2265 3328
rect 2122 3288 2126 3291
rect 2014 3282 2017 3288
rect 2182 3282 2185 3288
rect 2238 3282 2241 3288
rect 2074 3278 2078 3281
rect 2146 3278 2150 3281
rect 2078 3262 2081 3268
rect 2086 3262 2089 3278
rect 2110 3262 2113 3268
rect 2034 3258 2038 3261
rect 2058 3258 2062 3261
rect 2126 3252 2129 3268
rect 2254 3262 2257 3288
rect 2262 3262 2265 3278
rect 2138 3258 2142 3261
rect 2210 3258 2214 3261
rect 1962 3178 1966 3181
rect 2110 3162 2113 3168
rect 2134 3162 2137 3218
rect 2158 3182 2161 3258
rect 2198 3242 2201 3258
rect 2230 3252 2233 3258
rect 2222 3232 2225 3238
rect 2250 3228 2254 3231
rect 1902 3151 1905 3158
rect 1934 3152 1937 3158
rect 1970 3148 1974 3151
rect 2010 3148 2014 3151
rect 2030 3142 2033 3158
rect 2134 3152 2137 3158
rect 2050 3147 2054 3150
rect 2146 3148 2150 3151
rect 2166 3142 2169 3168
rect 2222 3152 2225 3158
rect 1978 3138 1982 3141
rect 2162 3138 2166 3141
rect 2118 3132 2121 3138
rect 2190 3132 2193 3138
rect 2230 3132 2233 3168
rect 2246 3152 2249 3168
rect 2270 3162 2273 3328
rect 2294 3302 2297 3328
rect 2278 3292 2281 3298
rect 2302 3292 2305 3328
rect 2326 3292 2329 3328
rect 2350 3292 2353 3328
rect 2406 3328 2418 3331
rect 2430 3328 2442 3331
rect 2470 3328 2474 3332
rect 2486 3328 2490 3332
rect 2502 3331 2506 3332
rect 2494 3328 2506 3331
rect 2526 3328 2530 3332
rect 2558 3328 2562 3332
rect 2574 3331 2578 3332
rect 2598 3331 2602 3332
rect 2574 3328 2585 3331
rect 2598 3328 2609 3331
rect 2406 3292 2409 3328
rect 2430 3292 2433 3328
rect 2470 3302 2473 3328
rect 2486 3292 2489 3328
rect 2494 3292 2497 3328
rect 2526 3302 2529 3328
rect 2558 3292 2561 3328
rect 2582 3292 2585 3328
rect 2606 3292 2609 3328
rect 2630 3328 2634 3332
rect 2646 3328 2650 3332
rect 2662 3328 2666 3332
rect 2678 3331 2682 3332
rect 2678 3328 2689 3331
rect 2630 3302 2633 3328
rect 2646 3292 2649 3328
rect 2662 3302 2665 3328
rect 2686 3292 2689 3328
rect 2766 3328 2770 3332
rect 2798 3328 2802 3332
rect 2814 3328 2818 3332
rect 2926 3328 2930 3332
rect 2942 3328 2946 3332
rect 2958 3328 2962 3332
rect 2974 3328 2978 3332
rect 2990 3331 2994 3332
rect 3014 3331 3018 3332
rect 2990 3328 3001 3331
rect 3014 3328 3025 3331
rect 2394 3288 2398 3291
rect 2474 3288 2478 3291
rect 2630 3282 2633 3288
rect 2666 3278 2670 3281
rect 2374 3272 2377 3278
rect 2306 3258 2310 3261
rect 2286 3242 2289 3258
rect 2334 3222 2337 3258
rect 2358 3222 2361 3258
rect 2398 3252 2401 3278
rect 2502 3272 2505 3278
rect 2454 3262 2457 3268
rect 2426 3258 2430 3261
rect 2506 3258 2510 3261
rect 2438 3192 2441 3238
rect 2446 3212 2449 3258
rect 2478 3172 2481 3258
rect 2518 3251 2521 3278
rect 2638 3272 2641 3278
rect 2694 3272 2697 3278
rect 2526 3262 2529 3268
rect 2518 3248 2526 3251
rect 2338 3158 2342 3161
rect 2474 3158 2478 3161
rect 2002 3128 2006 3131
rect 2130 3128 2134 3131
rect 2170 3128 2174 3131
rect 1886 3072 1889 3078
rect 1894 3021 1897 3098
rect 1998 3092 2001 3118
rect 2024 3103 2026 3107
rect 2030 3103 2033 3107
rect 2037 3103 2040 3107
rect 1954 3088 1958 3091
rect 1926 3072 1929 3078
rect 1990 3072 1993 3088
rect 2006 3082 2009 3088
rect 2046 3082 2049 3098
rect 2134 3092 2137 3108
rect 2142 3082 2145 3088
rect 2154 3078 2158 3081
rect 2062 3072 2065 3078
rect 2086 3072 2089 3078
rect 2094 3072 2097 3078
rect 2150 3072 2153 3078
rect 2010 3068 2014 3071
rect 2106 3068 2110 3071
rect 1902 3032 1905 3058
rect 1918 3052 1921 3068
rect 1894 3018 1905 3021
rect 1902 2992 1905 3018
rect 1838 2952 1841 2978
rect 1862 2962 1865 2968
rect 1830 2942 1833 2948
rect 1794 2928 1798 2931
rect 1806 2922 1809 2928
rect 1814 2901 1817 2918
rect 1838 2912 1841 2948
rect 1870 2942 1873 2978
rect 1886 2962 1889 2988
rect 1894 2962 1897 2968
rect 1926 2962 1929 3058
rect 1974 3042 1977 3068
rect 2070 3062 2073 3068
rect 2102 3062 2105 3068
rect 2126 3062 2129 3068
rect 1982 3052 1985 3058
rect 2014 3052 2017 3058
rect 1878 2942 1881 2948
rect 1850 2938 1854 2941
rect 1866 2928 1870 2931
rect 1814 2898 1822 2901
rect 1838 2892 1841 2898
rect 1870 2892 1873 2908
rect 1886 2882 1889 2958
rect 1950 2952 1953 3038
rect 1982 2962 1985 3028
rect 2046 2992 2049 3038
rect 2078 3032 2081 3058
rect 2102 2992 2105 3048
rect 2110 3032 2113 3058
rect 2118 3052 2121 3058
rect 2158 3032 2161 3068
rect 1990 2972 1993 2978
rect 2046 2962 2049 2978
rect 2062 2962 2065 2968
rect 2122 2958 2145 2961
rect 2154 2958 2158 2961
rect 1894 2942 1897 2948
rect 1918 2942 1921 2948
rect 2014 2942 2017 2948
rect 2038 2942 2041 2958
rect 1930 2938 1934 2941
rect 1986 2938 1990 2941
rect 2002 2938 2006 2941
rect 2046 2941 2049 2958
rect 2058 2948 2062 2951
rect 2046 2938 2054 2941
rect 1894 2892 1897 2918
rect 1918 2892 1921 2908
rect 1934 2902 1937 2918
rect 1850 2878 1854 2881
rect 1874 2878 1878 2881
rect 1650 2868 1654 2871
rect 1614 2842 1617 2848
rect 1638 2812 1641 2858
rect 1662 2842 1665 2848
rect 1590 2742 1593 2808
rect 1602 2758 1606 2761
rect 1630 2752 1633 2758
rect 1634 2738 1638 2741
rect 1582 2732 1585 2738
rect 1590 2682 1593 2738
rect 1642 2728 1646 2731
rect 1654 2722 1657 2728
rect 1606 2672 1609 2718
rect 1614 2712 1617 2718
rect 1594 2668 1598 2671
rect 1618 2668 1622 2671
rect 1550 2658 1558 2661
rect 1558 2652 1561 2658
rect 1574 2652 1577 2658
rect 1538 2648 1542 2651
rect 1582 2642 1585 2658
rect 1594 2648 1598 2651
rect 1478 2562 1481 2588
rect 1494 2561 1497 2618
rect 1512 2603 1514 2607
rect 1518 2603 1521 2607
rect 1525 2603 1528 2607
rect 1550 2592 1553 2608
rect 1558 2592 1561 2618
rect 1574 2592 1577 2598
rect 1490 2558 1497 2561
rect 1458 2548 1462 2551
rect 1438 2542 1441 2548
rect 1410 2528 1414 2531
rect 1426 2528 1430 2531
rect 1406 2482 1409 2488
rect 1414 2482 1417 2528
rect 1454 2522 1457 2538
rect 1470 2532 1473 2548
rect 1518 2532 1521 2548
rect 1526 2542 1529 2558
rect 1550 2552 1553 2588
rect 1582 2552 1585 2638
rect 1614 2612 1617 2658
rect 1590 2562 1593 2598
rect 1622 2552 1625 2648
rect 1538 2548 1542 2551
rect 1558 2542 1561 2548
rect 1546 2538 1550 2541
rect 1570 2538 1574 2541
rect 1446 2502 1449 2518
rect 1478 2512 1481 2518
rect 1450 2488 1454 2491
rect 1462 2472 1465 2478
rect 1378 2468 1385 2471
rect 1406 2468 1414 2471
rect 1266 2448 1273 2451
rect 1214 2402 1217 2418
rect 1246 2402 1249 2418
rect 1214 2362 1217 2368
rect 1234 2348 1238 2351
rect 1246 2342 1249 2348
rect 1254 2342 1257 2348
rect 1130 2338 1134 2341
rect 1142 2311 1145 2318
rect 1142 2308 1153 2311
rect 1142 2272 1145 2298
rect 1118 2242 1121 2248
rect 1126 2202 1129 2258
rect 1142 2252 1145 2258
rect 1150 2252 1153 2308
rect 1166 2282 1169 2328
rect 1174 2302 1177 2318
rect 1166 2262 1169 2278
rect 1174 2262 1177 2288
rect 1182 2272 1185 2278
rect 1190 2272 1193 2338
rect 1222 2312 1225 2318
rect 1150 2242 1153 2248
rect 1206 2242 1209 2248
rect 1214 2232 1217 2248
rect 1134 2162 1137 2228
rect 1190 2222 1193 2228
rect 1166 2202 1169 2218
rect 1166 2152 1169 2168
rect 1190 2152 1193 2158
rect 1198 2152 1201 2158
rect 1222 2152 1225 2298
rect 1230 2262 1233 2278
rect 1238 2272 1241 2298
rect 1246 2252 1249 2338
rect 1262 2291 1265 2398
rect 1270 2361 1273 2448
rect 1278 2382 1281 2418
rect 1286 2362 1289 2458
rect 1382 2452 1385 2458
rect 1270 2358 1278 2361
rect 1286 2342 1289 2358
rect 1254 2288 1265 2291
rect 1278 2292 1281 2318
rect 1286 2302 1289 2338
rect 1246 2242 1249 2248
rect 1254 2241 1257 2288
rect 1262 2272 1265 2278
rect 1270 2272 1273 2278
rect 1294 2272 1297 2448
rect 1326 2442 1329 2448
rect 1390 2442 1393 2458
rect 1302 2362 1305 2408
rect 1374 2402 1377 2418
rect 1398 2412 1401 2468
rect 1406 2462 1409 2468
rect 1430 2462 1433 2468
rect 1326 2392 1329 2398
rect 1338 2368 1342 2371
rect 1374 2362 1377 2378
rect 1350 2352 1353 2358
rect 1398 2352 1401 2358
rect 1338 2348 1342 2351
rect 1302 2342 1305 2348
rect 1406 2342 1409 2348
rect 1358 2332 1361 2338
rect 1322 2318 1326 2321
rect 1294 2262 1297 2268
rect 1278 2242 1281 2258
rect 1302 2251 1305 2318
rect 1342 2262 1345 2298
rect 1350 2272 1353 2278
rect 1382 2272 1385 2318
rect 1398 2272 1401 2288
rect 1298 2248 1305 2251
rect 1334 2252 1337 2258
rect 1254 2238 1265 2241
rect 1254 2222 1257 2228
rect 1230 2192 1233 2218
rect 1262 2162 1265 2238
rect 1350 2232 1353 2268
rect 1414 2262 1417 2458
rect 1462 2452 1465 2468
rect 1470 2462 1473 2498
rect 1494 2472 1497 2518
rect 1502 2462 1505 2498
rect 1558 2472 1561 2538
rect 1582 2492 1585 2548
rect 1606 2532 1609 2548
rect 1630 2541 1633 2708
rect 1646 2682 1649 2718
rect 1654 2682 1657 2718
rect 1662 2672 1665 2738
rect 1670 2722 1673 2858
rect 1702 2832 1705 2868
rect 1718 2852 1721 2858
rect 1698 2818 1702 2821
rect 1726 2812 1729 2868
rect 1782 2862 1785 2868
rect 1678 2732 1681 2808
rect 1694 2762 1697 2768
rect 1702 2742 1705 2758
rect 1642 2668 1646 2671
rect 1670 2662 1673 2678
rect 1678 2672 1681 2728
rect 1702 2691 1705 2738
rect 1710 2732 1713 2748
rect 1734 2732 1737 2858
rect 1754 2848 1758 2851
rect 1774 2851 1777 2858
rect 1770 2848 1777 2851
rect 1786 2848 1790 2851
rect 1806 2842 1809 2858
rect 1814 2852 1817 2868
rect 1822 2862 1825 2878
rect 1910 2871 1913 2878
rect 1910 2868 1921 2871
rect 1746 2838 1750 2841
rect 1806 2812 1809 2818
rect 1806 2762 1809 2768
rect 1822 2762 1825 2768
rect 1698 2688 1705 2691
rect 1694 2682 1697 2688
rect 1686 2672 1689 2678
rect 1718 2672 1721 2718
rect 1726 2692 1729 2728
rect 1726 2682 1729 2688
rect 1678 2662 1681 2668
rect 1694 2662 1697 2668
rect 1734 2662 1737 2728
rect 1742 2662 1745 2748
rect 1774 2722 1777 2738
rect 1782 2732 1785 2748
rect 1750 2682 1753 2718
rect 1782 2712 1785 2728
rect 1782 2672 1785 2678
rect 1762 2668 1766 2671
rect 1790 2662 1793 2758
rect 1798 2722 1801 2748
rect 1806 2732 1809 2738
rect 1806 2682 1809 2688
rect 1814 2662 1817 2718
rect 1830 2692 1833 2868
rect 1846 2862 1849 2868
rect 1854 2762 1857 2858
rect 1902 2852 1905 2858
rect 1902 2832 1905 2848
rect 1870 2752 1873 2768
rect 1882 2758 1886 2761
rect 1858 2748 1862 2751
rect 1902 2748 1910 2751
rect 1858 2738 1862 2741
rect 1894 2732 1897 2738
rect 1902 2722 1905 2748
rect 1918 2742 1921 2868
rect 1926 2862 1929 2868
rect 1950 2862 1953 2878
rect 1930 2848 1934 2851
rect 1946 2848 1950 2851
rect 1958 2822 1961 2938
rect 2070 2932 2073 2958
rect 2142 2952 2145 2958
rect 2082 2948 2086 2951
rect 2106 2948 2110 2951
rect 2166 2951 2169 3098
rect 2182 3082 2185 3118
rect 2186 3068 2190 3071
rect 2206 3062 2209 3128
rect 2230 3082 2233 3088
rect 2198 3052 2201 3058
rect 2174 2962 2177 2968
rect 2206 2962 2209 3028
rect 2214 3002 2217 3058
rect 2230 2982 2233 3048
rect 2238 3002 2241 3118
rect 2246 3092 2249 3148
rect 2270 3142 2273 3158
rect 2294 3152 2297 3158
rect 2326 3152 2329 3158
rect 2342 3142 2345 3148
rect 2306 3138 2310 3141
rect 2254 3132 2257 3138
rect 2262 3082 2265 3118
rect 2270 3102 2273 3138
rect 2290 3088 2294 3091
rect 2266 3078 2273 3081
rect 2270 3072 2273 3078
rect 2262 3042 2265 3068
rect 2286 3062 2289 3068
rect 2302 3051 2305 3118
rect 2358 3082 2361 3138
rect 2374 3112 2377 3147
rect 2390 3112 2393 3138
rect 2422 3092 2425 3158
rect 2486 3152 2489 3168
rect 2498 3158 2502 3161
rect 2526 3152 2529 3248
rect 2536 3203 2538 3207
rect 2542 3203 2545 3207
rect 2549 3203 2552 3207
rect 2454 3122 2457 3128
rect 2462 3102 2465 3128
rect 2470 3122 2473 3128
rect 2494 3092 2497 3128
rect 2510 3122 2513 3128
rect 2510 3102 2513 3118
rect 2518 3082 2521 3118
rect 2534 3092 2537 3138
rect 2558 3121 2561 3258
rect 2590 3252 2593 3258
rect 2614 3242 2617 3258
rect 2574 3142 2577 3147
rect 2550 3118 2561 3121
rect 2434 3078 2438 3081
rect 2538 3078 2542 3081
rect 2390 3072 2393 3078
rect 2446 3072 2449 3078
rect 2470 3072 2473 3078
rect 2458 3068 2462 3071
rect 2346 3058 2350 3061
rect 2290 3048 2305 3051
rect 2186 2958 2190 2961
rect 2206 2952 2209 2958
rect 2222 2952 2225 2958
rect 2166 2948 2174 2951
rect 2082 2938 2086 2941
rect 1990 2922 1993 2928
rect 2024 2903 2026 2907
rect 2030 2903 2033 2907
rect 2037 2903 2040 2907
rect 1966 2872 1969 2878
rect 1966 2852 1969 2858
rect 1974 2782 1977 2868
rect 1982 2862 1985 2878
rect 1994 2858 1998 2861
rect 2006 2832 2009 2868
rect 1926 2752 1929 2768
rect 1970 2758 1977 2761
rect 1974 2752 1977 2758
rect 1914 2738 1918 2741
rect 1838 2692 1841 2718
rect 1910 2691 1913 2738
rect 1902 2688 1913 2691
rect 1926 2692 1929 2718
rect 1966 2692 1969 2748
rect 1974 2732 1977 2738
rect 1822 2672 1825 2678
rect 1686 2658 1694 2661
rect 1654 2612 1657 2658
rect 1678 2562 1681 2598
rect 1646 2552 1649 2558
rect 1674 2548 1678 2551
rect 1630 2538 1638 2541
rect 1614 2532 1617 2538
rect 1590 2492 1593 2518
rect 1586 2478 1590 2481
rect 1422 2432 1425 2438
rect 1422 2392 1425 2408
rect 1394 2258 1398 2261
rect 1430 2261 1433 2378
rect 1454 2352 1457 2358
rect 1438 2292 1441 2348
rect 1462 2342 1465 2388
rect 1478 2351 1481 2368
rect 1486 2362 1489 2458
rect 1498 2448 1502 2451
rect 1522 2448 1526 2451
rect 1514 2438 1518 2441
rect 1512 2403 1514 2407
rect 1518 2403 1521 2407
rect 1525 2403 1528 2407
rect 1474 2348 1481 2351
rect 1454 2312 1457 2328
rect 1478 2282 1481 2348
rect 1498 2338 1502 2341
rect 1510 2282 1513 2388
rect 1526 2352 1529 2358
rect 1534 2352 1537 2468
rect 1566 2452 1569 2468
rect 1574 2462 1577 2478
rect 1598 2462 1601 2498
rect 1606 2481 1609 2518
rect 1622 2482 1625 2528
rect 1654 2522 1657 2538
rect 1634 2518 1641 2521
rect 1630 2492 1633 2508
rect 1606 2478 1614 2481
rect 1638 2472 1641 2518
rect 1662 2511 1665 2548
rect 1686 2542 1689 2658
rect 1722 2648 1726 2651
rect 1774 2642 1777 2658
rect 1710 2602 1713 2618
rect 1694 2552 1697 2558
rect 1702 2552 1705 2558
rect 1722 2548 1729 2551
rect 1738 2548 1742 2551
rect 1686 2532 1689 2538
rect 1654 2508 1665 2511
rect 1654 2502 1657 2508
rect 1662 2472 1665 2488
rect 1678 2482 1681 2488
rect 1686 2482 1689 2498
rect 1702 2482 1705 2548
rect 1726 2542 1729 2548
rect 1738 2538 1742 2541
rect 1610 2468 1614 2471
rect 1542 2392 1545 2448
rect 1554 2438 1558 2441
rect 1550 2342 1553 2408
rect 1562 2388 1566 2391
rect 1574 2372 1577 2458
rect 1586 2448 1590 2451
rect 1646 2402 1649 2458
rect 1654 2392 1657 2458
rect 1678 2442 1681 2448
rect 1686 2392 1689 2468
rect 1702 2412 1705 2478
rect 1602 2358 1606 2361
rect 1614 2352 1617 2358
rect 1662 2352 1665 2358
rect 1574 2342 1577 2348
rect 1654 2342 1657 2348
rect 1542 2338 1550 2341
rect 1610 2338 1614 2341
rect 1522 2328 1526 2331
rect 1542 2292 1545 2338
rect 1566 2292 1569 2328
rect 1590 2312 1593 2318
rect 1598 2302 1601 2338
rect 1634 2328 1638 2331
rect 1654 2302 1657 2328
rect 1450 2278 1454 2281
rect 1498 2278 1502 2281
rect 1470 2272 1473 2278
rect 1446 2262 1449 2268
rect 1478 2262 1481 2278
rect 1534 2272 1537 2278
rect 1542 2272 1545 2288
rect 1566 2282 1569 2288
rect 1590 2278 1614 2281
rect 1550 2262 1553 2278
rect 1574 2272 1577 2278
rect 1590 2272 1593 2278
rect 1630 2272 1633 2288
rect 1678 2272 1681 2328
rect 1562 2268 1566 2271
rect 1610 2268 1614 2271
rect 1650 2268 1654 2271
rect 1582 2262 1585 2268
rect 1430 2258 1438 2261
rect 1370 2248 1374 2251
rect 1278 2202 1281 2218
rect 1310 2162 1313 2188
rect 1326 2162 1329 2218
rect 1282 2158 1286 2161
rect 1254 2152 1257 2158
rect 1154 2148 1158 2151
rect 1282 2148 1286 2151
rect 998 2142 1001 2148
rect 1118 2142 1121 2148
rect 1334 2142 1337 2148
rect 1066 2138 1070 2141
rect 1166 2138 1174 2141
rect 982 2118 993 2121
rect 886 2061 889 2118
rect 910 2102 913 2118
rect 894 2078 913 2081
rect 922 2078 926 2081
rect 894 2072 897 2078
rect 910 2071 913 2078
rect 950 2072 953 2088
rect 910 2068 950 2071
rect 878 2058 889 2061
rect 902 2062 905 2068
rect 822 2048 830 2051
rect 762 1948 766 1951
rect 762 1938 766 1941
rect 750 1932 753 1938
rect 678 1882 681 1898
rect 650 1858 654 1861
rect 686 1861 689 1918
rect 694 1902 697 1928
rect 714 1868 718 1871
rect 678 1858 689 1861
rect 634 1758 641 1761
rect 638 1751 641 1758
rect 638 1748 646 1751
rect 610 1738 614 1741
rect 590 1722 593 1738
rect 598 1682 601 1688
rect 550 1678 561 1681
rect 526 1662 529 1668
rect 494 1648 502 1651
rect 390 1552 393 1608
rect 406 1602 409 1618
rect 480 1603 482 1607
rect 486 1603 489 1607
rect 493 1603 496 1607
rect 418 1568 422 1571
rect 398 1562 401 1568
rect 446 1562 449 1568
rect 470 1562 473 1568
rect 502 1561 505 1648
rect 530 1638 534 1641
rect 526 1562 529 1568
rect 502 1558 513 1561
rect 414 1542 417 1548
rect 450 1538 454 1541
rect 490 1538 494 1541
rect 374 1522 377 1528
rect 374 1462 377 1478
rect 382 1472 385 1518
rect 390 1472 393 1488
rect 414 1472 417 1538
rect 422 1532 425 1538
rect 502 1522 505 1548
rect 442 1518 446 1521
rect 450 1488 454 1491
rect 422 1472 425 1478
rect 398 1452 401 1458
rect 414 1452 417 1458
rect 374 1382 377 1418
rect 390 1362 393 1448
rect 398 1432 401 1448
rect 398 1362 401 1398
rect 354 1358 358 1361
rect 322 1348 326 1351
rect 322 1338 326 1341
rect 310 1332 313 1338
rect 318 1272 321 1298
rect 342 1292 345 1318
rect 350 1282 353 1318
rect 366 1292 369 1348
rect 414 1342 417 1438
rect 422 1362 425 1368
rect 374 1302 377 1338
rect 290 1268 294 1271
rect 250 1248 254 1251
rect 242 1238 246 1241
rect 174 1158 182 1161
rect 194 1148 198 1151
rect 142 1142 145 1148
rect 206 1142 209 1148
rect 214 1142 217 1238
rect 238 1182 241 1188
rect 222 1162 225 1168
rect 86 1092 89 1118
rect 26 1058 33 1061
rect 42 1078 46 1081
rect 74 1078 78 1081
rect 10 1048 14 1051
rect 6 962 9 968
rect 22 942 25 1058
rect 30 992 33 1038
rect 38 972 41 1078
rect 58 1068 62 1071
rect 94 1061 97 1138
rect 110 1132 113 1138
rect 134 1132 137 1138
rect 118 1102 121 1118
rect 90 1058 97 1061
rect 74 1048 78 1051
rect 86 1012 89 1058
rect 110 1052 113 1078
rect 138 1068 142 1071
rect 166 1071 169 1118
rect 174 1092 177 1108
rect 158 1068 169 1071
rect 182 1072 185 1138
rect 238 1072 241 1148
rect 254 1122 257 1128
rect 194 1068 198 1071
rect 118 1062 121 1068
rect 118 1042 121 1058
rect 134 1052 137 1068
rect 150 1062 153 1068
rect 146 1058 150 1061
rect 158 1051 161 1068
rect 170 1058 174 1061
rect 158 1048 166 1051
rect 86 962 89 968
rect 82 948 86 951
rect 70 942 73 948
rect 94 942 97 1038
rect 126 1032 129 1038
rect 126 992 129 1018
rect 102 962 105 968
rect 110 952 113 958
rect 114 948 121 951
rect 26 938 30 941
rect 86 938 94 941
rect 14 882 17 918
rect 38 892 41 928
rect 46 912 49 928
rect 10 868 14 871
rect 30 851 33 878
rect 62 872 65 878
rect 42 858 49 861
rect 30 848 38 851
rect 46 812 49 858
rect 70 861 73 938
rect 86 872 89 938
rect 118 932 121 948
rect 134 942 137 1008
rect 150 962 153 1048
rect 174 1042 177 1048
rect 158 962 161 968
rect 182 952 185 1068
rect 238 1062 241 1068
rect 190 972 193 1018
rect 198 961 201 1058
rect 206 1042 209 1058
rect 254 1052 257 1118
rect 262 1092 265 1198
rect 270 1182 273 1258
rect 302 1252 305 1268
rect 318 1262 321 1268
rect 290 1248 294 1251
rect 318 1242 321 1258
rect 334 1252 337 1278
rect 318 1212 321 1218
rect 290 1168 294 1171
rect 310 1152 313 1208
rect 318 1162 321 1178
rect 274 1148 278 1151
rect 314 1148 318 1151
rect 302 1141 305 1148
rect 334 1142 337 1238
rect 342 1192 345 1268
rect 350 1262 353 1268
rect 358 1162 361 1278
rect 382 1272 385 1318
rect 366 1252 369 1268
rect 374 1252 377 1258
rect 302 1138 313 1141
rect 234 968 238 971
rect 270 962 273 1118
rect 310 1072 313 1138
rect 290 1068 294 1071
rect 298 1058 302 1061
rect 278 1042 281 1058
rect 286 972 289 1058
rect 318 1052 321 1118
rect 334 1062 337 1138
rect 342 1082 345 1148
rect 342 1072 345 1078
rect 350 1062 353 1068
rect 358 1051 361 1118
rect 374 1102 377 1148
rect 390 1142 393 1298
rect 398 1282 401 1318
rect 414 1272 417 1338
rect 398 1262 401 1268
rect 402 1248 406 1251
rect 398 1182 401 1188
rect 414 1171 417 1268
rect 422 1262 425 1278
rect 430 1272 433 1448
rect 446 1372 449 1458
rect 454 1432 457 1468
rect 462 1462 465 1468
rect 470 1451 473 1518
rect 490 1468 494 1471
rect 466 1448 473 1451
rect 478 1442 481 1458
rect 480 1403 482 1407
rect 486 1403 489 1407
rect 493 1403 496 1407
rect 486 1362 489 1378
rect 466 1358 470 1361
rect 438 1352 441 1358
rect 458 1348 462 1351
rect 450 1338 454 1341
rect 438 1332 441 1338
rect 442 1328 449 1331
rect 446 1322 449 1328
rect 486 1292 489 1318
rect 438 1272 441 1278
rect 446 1272 449 1278
rect 430 1262 433 1268
rect 454 1262 457 1288
rect 494 1272 497 1388
rect 494 1262 497 1268
rect 502 1262 505 1518
rect 510 1462 513 1558
rect 542 1552 545 1598
rect 550 1552 553 1668
rect 558 1662 561 1678
rect 538 1538 542 1541
rect 518 1462 521 1518
rect 558 1472 561 1598
rect 566 1572 569 1658
rect 574 1652 577 1678
rect 582 1662 585 1668
rect 598 1662 601 1668
rect 614 1662 617 1718
rect 622 1672 625 1748
rect 642 1738 646 1741
rect 654 1731 657 1818
rect 662 1752 665 1758
rect 670 1751 673 1818
rect 678 1761 681 1858
rect 690 1848 694 1851
rect 726 1851 729 1918
rect 742 1912 745 1918
rect 774 1912 777 1938
rect 746 1868 750 1871
rect 766 1862 769 1868
rect 798 1862 801 1878
rect 814 1862 817 2018
rect 822 1942 825 1958
rect 838 1941 841 2058
rect 846 1952 849 2038
rect 854 1942 857 1948
rect 838 1938 846 1941
rect 822 1882 825 1918
rect 862 1912 865 2018
rect 878 1962 881 2058
rect 942 2052 945 2058
rect 922 2048 926 2051
rect 886 2042 889 2048
rect 886 1962 889 2038
rect 910 1982 913 2018
rect 926 1952 929 1968
rect 942 1952 945 2018
rect 950 1992 953 2058
rect 958 2052 961 2118
rect 982 2081 985 2118
rect 992 2103 994 2107
rect 998 2103 1001 2107
rect 1005 2103 1008 2107
rect 974 2078 985 2081
rect 974 2062 977 2078
rect 1002 2068 1006 2071
rect 982 2062 985 2068
rect 1014 2051 1017 2118
rect 1006 2048 1017 2051
rect 1030 2052 1033 2078
rect 1038 2072 1041 2088
rect 1046 2072 1049 2138
rect 1054 2082 1057 2118
rect 1070 2112 1073 2138
rect 1094 2132 1097 2138
rect 1110 2132 1113 2138
rect 1106 2118 1110 2121
rect 1050 2058 1054 2061
rect 1070 2052 1073 2088
rect 1006 2032 1009 2048
rect 1014 2032 1017 2038
rect 1046 1992 1049 2018
rect 958 1962 961 1978
rect 1022 1972 1025 1978
rect 966 1962 969 1968
rect 1038 1962 1041 1968
rect 1062 1962 1065 2038
rect 922 1948 926 1951
rect 1018 1948 1022 1951
rect 906 1938 910 1941
rect 870 1902 873 1938
rect 822 1862 825 1878
rect 834 1868 838 1871
rect 866 1868 870 1871
rect 778 1858 782 1861
rect 842 1858 846 1861
rect 758 1852 761 1858
rect 722 1848 729 1851
rect 738 1848 742 1851
rect 678 1758 686 1761
rect 670 1748 678 1751
rect 646 1728 657 1731
rect 646 1722 649 1728
rect 630 1682 633 1718
rect 678 1712 681 1718
rect 646 1672 649 1688
rect 654 1682 657 1708
rect 686 1691 689 1758
rect 702 1752 705 1818
rect 718 1772 721 1778
rect 710 1752 713 1768
rect 734 1762 737 1838
rect 738 1748 742 1751
rect 698 1738 702 1741
rect 714 1738 718 1741
rect 678 1688 689 1691
rect 678 1682 681 1688
rect 662 1672 665 1678
rect 686 1672 689 1678
rect 634 1668 638 1671
rect 626 1658 630 1661
rect 606 1602 609 1618
rect 598 1571 601 1588
rect 598 1568 609 1571
rect 566 1558 593 1561
rect 566 1552 569 1558
rect 590 1552 593 1558
rect 598 1552 601 1558
rect 578 1548 582 1551
rect 606 1551 609 1568
rect 630 1562 633 1598
rect 670 1591 673 1618
rect 662 1588 673 1591
rect 662 1552 665 1588
rect 606 1548 614 1551
rect 626 1548 630 1551
rect 578 1538 585 1541
rect 570 1528 574 1531
rect 582 1502 585 1538
rect 606 1532 609 1538
rect 598 1482 601 1518
rect 614 1472 617 1548
rect 654 1542 657 1548
rect 602 1468 606 1471
rect 538 1458 542 1461
rect 562 1458 566 1461
rect 622 1461 625 1538
rect 638 1512 641 1518
rect 618 1458 625 1461
rect 550 1452 553 1458
rect 590 1442 593 1458
rect 598 1452 601 1458
rect 638 1452 641 1498
rect 670 1492 673 1578
rect 650 1468 654 1471
rect 662 1462 665 1468
rect 618 1438 622 1441
rect 510 1392 513 1418
rect 526 1352 529 1368
rect 534 1362 537 1418
rect 582 1412 585 1418
rect 606 1372 609 1378
rect 570 1358 574 1361
rect 558 1352 561 1358
rect 606 1352 609 1358
rect 506 1258 513 1261
rect 454 1252 457 1258
rect 482 1248 486 1251
rect 422 1242 425 1248
rect 414 1168 425 1171
rect 414 1152 417 1158
rect 398 1142 401 1148
rect 422 1142 425 1168
rect 446 1162 449 1188
rect 442 1148 446 1151
rect 434 1118 438 1121
rect 454 1112 457 1238
rect 470 1152 473 1208
rect 480 1203 482 1207
rect 486 1203 489 1207
rect 493 1203 496 1207
rect 502 1192 505 1198
rect 510 1162 513 1258
rect 518 1222 521 1338
rect 526 1272 529 1348
rect 534 1342 537 1348
rect 586 1338 590 1341
rect 626 1338 630 1341
rect 550 1312 553 1318
rect 558 1272 561 1338
rect 558 1262 561 1268
rect 566 1262 569 1268
rect 534 1152 537 1218
rect 550 1192 553 1258
rect 582 1252 585 1318
rect 598 1272 601 1328
rect 638 1292 641 1388
rect 646 1362 649 1438
rect 646 1322 649 1338
rect 630 1272 633 1278
rect 594 1268 598 1271
rect 618 1268 622 1271
rect 606 1262 609 1268
rect 646 1262 649 1318
rect 654 1262 657 1378
rect 662 1341 665 1458
rect 678 1452 681 1598
rect 686 1532 689 1668
rect 694 1662 697 1718
rect 710 1652 713 1678
rect 742 1672 745 1708
rect 738 1658 742 1661
rect 750 1652 753 1668
rect 758 1662 761 1798
rect 766 1752 769 1858
rect 786 1848 790 1851
rect 774 1792 777 1818
rect 798 1802 801 1858
rect 798 1762 801 1788
rect 806 1762 809 1808
rect 814 1792 817 1818
rect 822 1762 825 1768
rect 766 1742 769 1748
rect 774 1742 777 1748
rect 790 1671 793 1728
rect 798 1702 801 1718
rect 806 1682 809 1718
rect 790 1668 798 1671
rect 806 1662 809 1668
rect 782 1652 785 1658
rect 718 1642 721 1648
rect 734 1632 737 1638
rect 758 1622 761 1628
rect 694 1602 697 1618
rect 722 1578 726 1581
rect 774 1562 777 1568
rect 726 1552 729 1558
rect 790 1552 793 1618
rect 798 1582 801 1658
rect 814 1612 817 1708
rect 822 1692 825 1738
rect 846 1732 849 1738
rect 854 1702 857 1718
rect 850 1668 854 1671
rect 834 1658 838 1661
rect 826 1648 830 1651
rect 846 1642 849 1658
rect 862 1652 865 1858
rect 878 1752 881 1908
rect 886 1872 889 1928
rect 910 1881 913 1918
rect 934 1902 937 1938
rect 942 1932 945 1938
rect 906 1878 913 1881
rect 938 1868 942 1871
rect 886 1742 889 1868
rect 918 1862 921 1868
rect 910 1762 913 1818
rect 918 1782 921 1858
rect 926 1802 929 1858
rect 918 1762 921 1768
rect 934 1742 937 1828
rect 950 1822 953 1918
rect 966 1882 969 1948
rect 1030 1942 1033 1958
rect 1070 1952 1073 2048
rect 1078 2042 1081 2118
rect 1086 2072 1089 2118
rect 1142 2092 1145 2118
rect 1102 2082 1105 2088
rect 1110 2052 1113 2068
rect 1118 2062 1121 2078
rect 1166 2072 1169 2138
rect 1078 1952 1081 2028
rect 1094 2002 1097 2018
rect 1102 1972 1105 1978
rect 1126 1962 1129 1968
rect 1086 1942 1089 1958
rect 978 1938 982 1941
rect 1098 1938 1102 1941
rect 974 1902 977 1928
rect 992 1903 994 1907
rect 998 1903 1001 1907
rect 1005 1903 1008 1907
rect 982 1852 985 1878
rect 994 1868 998 1871
rect 962 1848 966 1851
rect 958 1762 961 1808
rect 966 1782 969 1848
rect 974 1761 977 1818
rect 990 1772 993 1818
rect 1014 1792 1017 1868
rect 1030 1852 1033 1858
rect 1014 1762 1017 1788
rect 1030 1762 1033 1768
rect 1038 1762 1041 1858
rect 1046 1852 1049 1918
rect 1054 1882 1057 1938
rect 1062 1882 1065 1918
rect 1086 1872 1089 1878
rect 1110 1862 1113 1888
rect 1054 1762 1057 1778
rect 974 1758 982 1761
rect 982 1742 985 1758
rect 1014 1752 1017 1758
rect 874 1738 878 1741
rect 1034 1738 1038 1741
rect 878 1722 881 1738
rect 934 1732 937 1738
rect 942 1732 945 1738
rect 958 1732 961 1738
rect 922 1728 929 1731
rect 910 1712 913 1718
rect 886 1682 889 1708
rect 898 1688 902 1691
rect 874 1668 878 1671
rect 910 1671 913 1698
rect 906 1668 913 1671
rect 798 1558 806 1561
rect 798 1552 801 1558
rect 814 1551 817 1608
rect 830 1562 833 1608
rect 806 1548 817 1551
rect 694 1542 697 1548
rect 710 1532 713 1538
rect 686 1522 689 1528
rect 694 1512 697 1528
rect 706 1518 710 1521
rect 702 1482 705 1488
rect 678 1361 681 1448
rect 686 1371 689 1458
rect 686 1368 697 1371
rect 694 1362 697 1368
rect 674 1358 681 1361
rect 686 1352 689 1358
rect 702 1352 705 1358
rect 662 1338 670 1341
rect 662 1322 665 1338
rect 662 1272 665 1298
rect 590 1252 593 1258
rect 614 1241 617 1258
rect 638 1252 641 1258
rect 602 1238 617 1241
rect 646 1232 649 1258
rect 566 1192 569 1218
rect 582 1162 585 1208
rect 554 1158 558 1161
rect 614 1152 617 1228
rect 462 1132 465 1138
rect 430 1092 433 1098
rect 502 1092 505 1108
rect 518 1102 521 1148
rect 530 1138 534 1141
rect 402 1088 406 1091
rect 462 1072 465 1078
rect 370 1068 374 1071
rect 466 1068 470 1071
rect 386 1058 390 1061
rect 358 1048 366 1051
rect 374 1051 377 1058
rect 406 1052 409 1068
rect 422 1062 425 1068
rect 454 1062 457 1068
rect 442 1058 446 1061
rect 374 1048 398 1051
rect 346 1038 350 1041
rect 302 982 305 988
rect 310 962 313 968
rect 198 958 206 961
rect 186 938 190 941
rect 82 868 86 871
rect 94 862 97 868
rect 66 858 73 861
rect 62 852 65 858
rect 54 842 57 848
rect 70 842 73 848
rect 54 792 57 828
rect 78 752 81 858
rect 110 852 113 868
rect 134 862 137 938
rect 166 932 169 938
rect 186 928 190 931
rect 142 892 145 908
rect 122 848 126 851
rect 150 851 153 918
rect 162 858 166 861
rect 146 848 153 851
rect 86 842 89 848
rect 94 762 97 838
rect 14 682 17 718
rect 30 712 33 748
rect 42 738 46 741
rect 66 738 70 741
rect 42 728 46 731
rect 66 728 70 731
rect 14 662 17 668
rect 22 592 25 698
rect 38 672 41 678
rect 10 548 14 551
rect 22 472 25 518
rect 30 492 33 658
rect 54 652 57 728
rect 70 672 73 678
rect 78 672 81 748
rect 110 742 113 848
rect 122 838 126 841
rect 174 832 177 918
rect 182 852 185 878
rect 198 872 201 958
rect 326 952 329 1008
rect 358 962 361 978
rect 274 948 278 951
rect 222 942 225 948
rect 246 942 249 948
rect 206 872 209 928
rect 214 902 217 918
rect 222 872 225 938
rect 230 872 233 928
rect 246 872 249 938
rect 254 932 257 948
rect 286 932 289 948
rect 334 942 337 948
rect 354 938 358 941
rect 270 922 273 928
rect 294 922 297 928
rect 286 882 289 888
rect 254 872 257 878
rect 206 862 209 868
rect 214 862 217 868
rect 234 858 238 861
rect 126 792 129 808
rect 150 792 153 798
rect 174 792 177 828
rect 182 792 185 848
rect 190 842 193 848
rect 198 792 201 858
rect 206 772 209 858
rect 214 848 222 851
rect 294 851 297 898
rect 310 892 313 918
rect 318 872 321 918
rect 326 882 329 938
rect 346 888 350 891
rect 366 882 369 938
rect 374 892 377 1028
rect 382 962 385 988
rect 390 942 393 948
rect 398 932 401 948
rect 326 862 329 878
rect 366 872 369 878
rect 306 858 310 861
rect 294 848 310 851
rect 214 792 217 848
rect 258 838 262 841
rect 238 792 241 818
rect 270 802 273 848
rect 334 822 337 868
rect 342 852 345 858
rect 334 782 337 818
rect 226 758 230 761
rect 126 738 134 741
rect 86 732 89 738
rect 94 672 97 738
rect 118 692 121 718
rect 78 662 81 668
rect 58 648 62 651
rect 86 651 89 668
rect 94 662 97 668
rect 78 648 89 651
rect 110 652 113 678
rect 126 671 129 738
rect 142 722 145 728
rect 158 692 161 758
rect 174 732 177 748
rect 246 742 249 768
rect 262 762 265 768
rect 318 762 321 768
rect 350 762 353 818
rect 358 812 361 858
rect 382 851 385 918
rect 406 882 409 938
rect 414 892 417 958
rect 422 952 425 1058
rect 446 992 449 1038
rect 470 992 473 1058
rect 478 1052 481 1088
rect 514 1058 518 1061
rect 526 1042 529 1068
rect 534 1052 537 1098
rect 480 1003 482 1007
rect 486 1003 489 1007
rect 493 1003 496 1007
rect 510 992 513 1038
rect 422 942 425 948
rect 398 872 401 878
rect 422 872 425 908
rect 430 902 433 948
rect 438 872 441 968
rect 454 952 457 988
rect 526 952 529 1008
rect 542 962 545 1118
rect 558 1092 561 1148
rect 606 1142 609 1148
rect 566 1072 569 1118
rect 550 1062 553 1068
rect 574 1062 577 1128
rect 590 1102 593 1118
rect 586 1068 590 1071
rect 606 1062 609 1138
rect 622 1082 625 1118
rect 618 1068 622 1071
rect 578 1058 582 1061
rect 610 1058 614 1061
rect 582 1048 590 1051
rect 582 1042 585 1048
rect 590 992 593 1038
rect 550 952 553 958
rect 526 942 529 948
rect 482 928 486 931
rect 478 892 481 898
rect 458 878 462 881
rect 482 878 486 881
rect 502 872 505 928
rect 518 882 521 938
rect 534 892 537 948
rect 542 932 545 938
rect 550 892 553 938
rect 558 902 561 938
rect 566 932 569 948
rect 574 942 577 958
rect 606 952 609 1018
rect 614 932 617 1058
rect 630 1031 633 1188
rect 654 1182 657 1258
rect 670 1252 673 1318
rect 686 1271 689 1348
rect 710 1342 713 1468
rect 718 1442 721 1538
rect 718 1352 721 1438
rect 726 1432 729 1548
rect 750 1542 753 1548
rect 758 1512 761 1538
rect 798 1482 801 1548
rect 806 1542 809 1548
rect 818 1538 822 1541
rect 738 1468 742 1471
rect 750 1462 753 1478
rect 766 1462 769 1468
rect 762 1448 766 1451
rect 774 1442 777 1468
rect 794 1448 798 1451
rect 806 1441 809 1538
rect 822 1502 825 1518
rect 822 1462 825 1488
rect 830 1462 833 1538
rect 838 1532 841 1568
rect 838 1492 841 1498
rect 846 1482 849 1608
rect 862 1572 865 1648
rect 882 1638 886 1641
rect 882 1578 897 1581
rect 894 1572 897 1578
rect 870 1542 873 1548
rect 862 1511 865 1518
rect 858 1508 865 1511
rect 870 1472 873 1528
rect 878 1512 881 1568
rect 886 1562 889 1568
rect 890 1558 897 1561
rect 894 1532 897 1558
rect 870 1462 873 1468
rect 894 1452 897 1478
rect 902 1462 905 1658
rect 918 1651 921 1718
rect 926 1712 929 1728
rect 930 1688 934 1691
rect 958 1672 961 1718
rect 966 1712 969 1738
rect 1058 1728 1062 1731
rect 930 1668 934 1671
rect 966 1662 969 1668
rect 918 1648 926 1651
rect 938 1648 942 1651
rect 910 1562 913 1568
rect 918 1561 921 1578
rect 930 1568 934 1571
rect 918 1558 929 1561
rect 926 1552 929 1558
rect 950 1552 953 1558
rect 914 1548 918 1551
rect 938 1548 942 1551
rect 926 1512 929 1548
rect 934 1532 937 1538
rect 958 1522 961 1528
rect 966 1511 969 1538
rect 974 1531 977 1658
rect 982 1652 985 1718
rect 992 1703 994 1707
rect 998 1703 1001 1707
rect 1005 1703 1008 1707
rect 1030 1702 1033 1718
rect 1014 1662 1017 1688
rect 1038 1662 1041 1668
rect 1054 1662 1057 1678
rect 1070 1671 1073 1838
rect 1078 1752 1081 1758
rect 1086 1742 1089 1778
rect 1094 1762 1097 1768
rect 1086 1712 1089 1738
rect 1102 1712 1105 1858
rect 1118 1792 1121 1868
rect 1134 1862 1137 2058
rect 1142 2052 1145 2068
rect 1166 2052 1169 2068
rect 1174 2062 1177 2078
rect 1190 2052 1193 2118
rect 1222 2092 1225 2138
rect 1246 2122 1249 2138
rect 1262 2102 1265 2118
rect 1278 2112 1281 2138
rect 1302 2132 1305 2138
rect 1326 2132 1329 2138
rect 1314 2118 1318 2121
rect 1142 1942 1145 2048
rect 1198 2042 1201 2048
rect 1174 1982 1177 2018
rect 1166 1952 1169 1958
rect 1190 1952 1193 1978
rect 1206 1952 1209 2088
rect 1214 2062 1217 2088
rect 1222 2072 1225 2088
rect 1178 1948 1182 1951
rect 1194 1938 1198 1941
rect 1206 1932 1209 1938
rect 1214 1912 1217 2018
rect 1222 1992 1225 2058
rect 1230 2052 1233 2098
rect 1286 2072 1289 2088
rect 1302 2072 1305 2108
rect 1326 2092 1329 2128
rect 1334 2072 1337 2088
rect 1342 2082 1345 2188
rect 1374 2162 1377 2198
rect 1382 2182 1385 2258
rect 1354 2158 1358 2161
rect 1398 2152 1401 2258
rect 1414 2252 1417 2258
rect 1438 2252 1441 2258
rect 1410 2158 1414 2161
rect 1314 2068 1318 2071
rect 1246 2052 1249 2058
rect 1262 2002 1265 2068
rect 1278 2052 1281 2068
rect 1302 2052 1305 2068
rect 1326 2062 1329 2068
rect 1270 1992 1273 2018
rect 1238 1962 1241 1968
rect 1270 1952 1273 1978
rect 1286 1962 1289 1988
rect 1350 1962 1353 2118
rect 1358 2092 1361 2138
rect 1366 2062 1369 2088
rect 1374 2051 1377 2118
rect 1382 2092 1385 2138
rect 1390 2062 1393 2088
rect 1398 2062 1401 2078
rect 1398 2052 1401 2058
rect 1374 2048 1382 2051
rect 1406 2032 1409 2118
rect 1422 2072 1425 2218
rect 1438 2152 1441 2238
rect 1446 2162 1449 2258
rect 1454 2151 1457 2258
rect 1598 2252 1601 2258
rect 1450 2148 1457 2151
rect 1470 2152 1473 2248
rect 1558 2242 1561 2248
rect 1486 2152 1489 2198
rect 1430 2092 1433 2138
rect 1502 2132 1505 2228
rect 1512 2203 1514 2207
rect 1518 2203 1521 2207
rect 1525 2203 1528 2207
rect 1514 2178 1518 2181
rect 1534 2172 1537 2178
rect 1522 2148 1534 2151
rect 1438 2092 1441 2098
rect 1422 2062 1425 2068
rect 1446 2062 1449 2078
rect 1454 2072 1457 2088
rect 1462 2062 1465 2118
rect 1486 2072 1489 2088
rect 1502 2062 1505 2128
rect 1510 2122 1513 2128
rect 1414 2042 1417 2048
rect 1502 2042 1505 2048
rect 1510 2042 1513 2118
rect 1550 2102 1553 2158
rect 1558 2152 1561 2178
rect 1606 2171 1609 2258
rect 1614 2182 1617 2218
rect 1598 2168 1609 2171
rect 1598 2162 1601 2168
rect 1610 2158 1638 2161
rect 1646 2152 1649 2258
rect 1686 2252 1689 2388
rect 1698 2348 1702 2351
rect 1710 2342 1713 2528
rect 1718 2512 1721 2518
rect 1734 2492 1737 2518
rect 1750 2492 1753 2618
rect 1790 2582 1793 2658
rect 1838 2622 1841 2678
rect 1894 2672 1897 2678
rect 1890 2668 1894 2671
rect 1870 2662 1873 2668
rect 1902 2662 1905 2688
rect 1914 2678 1918 2681
rect 1966 2671 1969 2678
rect 1962 2668 1969 2671
rect 1918 2662 1921 2668
rect 1942 2662 1945 2668
rect 1854 2652 1857 2658
rect 1902 2652 1905 2658
rect 1882 2648 1886 2651
rect 1846 2612 1849 2648
rect 1838 2598 1846 2601
rect 1838 2592 1841 2598
rect 1818 2588 1822 2591
rect 1770 2558 1777 2561
rect 1758 2552 1761 2558
rect 1822 2542 1825 2578
rect 1886 2562 1889 2618
rect 1858 2558 1881 2561
rect 1878 2552 1881 2558
rect 1894 2552 1897 2558
rect 1958 2552 1961 2558
rect 1858 2548 1862 2551
rect 1930 2548 1934 2551
rect 1830 2542 1833 2548
rect 1838 2542 1841 2548
rect 1786 2538 1790 2541
rect 1866 2538 1870 2541
rect 1718 2452 1721 2458
rect 1742 2452 1745 2478
rect 1766 2462 1769 2538
rect 1774 2501 1777 2518
rect 1782 2501 1785 2508
rect 1774 2498 1785 2501
rect 1774 2472 1777 2488
rect 1782 2462 1785 2498
rect 1790 2492 1793 2498
rect 1822 2482 1825 2488
rect 1830 2482 1833 2538
rect 1886 2532 1889 2538
rect 1910 2532 1913 2538
rect 1926 2522 1929 2528
rect 1854 2492 1857 2518
rect 1766 2452 1769 2458
rect 1798 2452 1801 2458
rect 1750 2422 1753 2448
rect 1770 2438 1774 2441
rect 1806 2422 1809 2478
rect 1826 2468 1830 2471
rect 1818 2448 1822 2451
rect 1838 2422 1841 2458
rect 1806 2392 1809 2418
rect 1854 2392 1857 2448
rect 1862 2422 1865 2478
rect 1878 2462 1881 2468
rect 1890 2418 1894 2421
rect 1902 2412 1905 2478
rect 1910 2452 1913 2468
rect 1926 2462 1929 2508
rect 1934 2482 1937 2538
rect 1942 2522 1945 2538
rect 1950 2501 1953 2548
rect 1966 2542 1969 2668
rect 1974 2592 1977 2708
rect 1982 2692 1985 2828
rect 1998 2772 2001 2818
rect 1990 2722 1993 2738
rect 2006 2722 2009 2728
rect 2006 2682 2009 2688
rect 1982 2532 1985 2538
rect 1946 2498 1953 2501
rect 1990 2502 1993 2538
rect 1942 2482 1945 2498
rect 1998 2492 2001 2608
rect 2006 2602 2009 2658
rect 2014 2642 2017 2858
rect 2022 2792 2025 2808
rect 2038 2782 2041 2868
rect 2054 2852 2057 2868
rect 2062 2862 2065 2918
rect 2070 2862 2073 2928
rect 2094 2922 2097 2938
rect 2126 2922 2129 2948
rect 2134 2942 2137 2948
rect 2182 2942 2185 2948
rect 2102 2872 2105 2898
rect 2118 2872 2121 2878
rect 2070 2841 2073 2848
rect 2058 2838 2073 2841
rect 2094 2832 2097 2868
rect 2118 2852 2121 2858
rect 2086 2762 2089 2818
rect 2114 2768 2118 2771
rect 2038 2732 2041 2738
rect 2024 2703 2026 2707
rect 2030 2703 2033 2707
rect 2037 2703 2040 2707
rect 2046 2692 2049 2758
rect 2054 2752 2057 2758
rect 2062 2682 2065 2748
rect 2110 2742 2113 2748
rect 2118 2742 2121 2748
rect 2074 2738 2078 2741
rect 2082 2728 2086 2731
rect 2134 2731 2137 2938
rect 2150 2912 2153 2928
rect 2150 2882 2153 2888
rect 2162 2868 2166 2871
rect 2162 2828 2166 2831
rect 2142 2742 2145 2828
rect 2174 2802 2177 2848
rect 2190 2832 2193 2918
rect 2198 2882 2201 2948
rect 2238 2942 2241 2978
rect 2214 2882 2217 2938
rect 2198 2872 2201 2878
rect 2206 2872 2209 2878
rect 2222 2872 2225 2938
rect 2230 2902 2233 2918
rect 2206 2852 2209 2868
rect 2218 2858 2222 2861
rect 2230 2852 2233 2898
rect 2238 2892 2241 2938
rect 2254 2931 2257 3018
rect 2278 2962 2281 3018
rect 2302 2962 2305 3038
rect 2330 2958 2334 2961
rect 2270 2942 2273 2948
rect 2278 2942 2281 2958
rect 2314 2938 2318 2941
rect 2250 2928 2257 2931
rect 2278 2932 2281 2938
rect 2326 2932 2329 2948
rect 2366 2942 2369 2947
rect 2374 2942 2377 3068
rect 2406 3062 2409 3068
rect 2486 3062 2489 3068
rect 2494 3062 2497 3068
rect 2422 3052 2425 3058
rect 2454 3052 2457 3058
rect 2502 3052 2505 3058
rect 2482 3048 2486 3051
rect 2430 3042 2433 3048
rect 2430 2992 2433 2998
rect 2438 2982 2441 3008
rect 2438 2932 2441 2938
rect 2254 2901 2257 2918
rect 2286 2902 2289 2918
rect 2254 2898 2265 2901
rect 2250 2888 2254 2891
rect 2250 2868 2254 2871
rect 2238 2862 2241 2868
rect 2190 2772 2193 2818
rect 2166 2762 2169 2768
rect 2182 2752 2185 2758
rect 2190 2742 2193 2748
rect 2198 2742 2201 2838
rect 2222 2762 2225 2798
rect 2246 2782 2249 2798
rect 2214 2752 2217 2758
rect 2234 2748 2238 2751
rect 2222 2742 2225 2748
rect 2246 2742 2249 2778
rect 2262 2772 2265 2898
rect 2286 2872 2289 2878
rect 2302 2862 2305 2888
rect 2274 2858 2278 2861
rect 2290 2858 2294 2861
rect 2274 2848 2278 2851
rect 2270 2782 2273 2848
rect 2302 2792 2305 2818
rect 2198 2732 2201 2738
rect 2254 2732 2257 2768
rect 2262 2752 2265 2758
rect 2270 2742 2273 2778
rect 2282 2758 2286 2761
rect 2278 2742 2281 2748
rect 2134 2728 2145 2731
rect 2178 2728 2182 2731
rect 2110 2682 2113 2728
rect 2126 2722 2129 2728
rect 2130 2718 2137 2721
rect 2134 2682 2137 2718
rect 2142 2692 2145 2728
rect 2166 2682 2169 2718
rect 2222 2702 2225 2718
rect 2238 2692 2241 2708
rect 2254 2682 2257 2688
rect 2066 2678 2070 2681
rect 2210 2678 2214 2681
rect 2242 2678 2246 2681
rect 2286 2681 2289 2758
rect 2298 2748 2302 2751
rect 2282 2678 2289 2681
rect 2302 2692 2305 2748
rect 2302 2682 2305 2688
rect 2098 2668 2102 2671
rect 2114 2668 2118 2671
rect 2022 2652 2025 2658
rect 2062 2642 2065 2668
rect 2094 2662 2097 2668
rect 2126 2662 2129 2678
rect 2158 2672 2161 2678
rect 2194 2668 2198 2671
rect 2218 2668 2222 2671
rect 2150 2662 2153 2668
rect 2158 2662 2161 2668
rect 2106 2658 2110 2661
rect 2006 2552 2009 2558
rect 2014 2552 2017 2568
rect 2034 2548 2038 2551
rect 2042 2538 2046 2541
rect 2014 2532 2017 2538
rect 2026 2528 2030 2531
rect 2024 2503 2026 2507
rect 2030 2503 2033 2507
rect 2037 2503 2040 2507
rect 1962 2488 1966 2491
rect 1990 2482 1993 2488
rect 2046 2482 2049 2528
rect 2054 2522 2057 2578
rect 2102 2562 2105 2578
rect 2094 2558 2102 2561
rect 2094 2542 2097 2558
rect 2126 2542 2129 2548
rect 2086 2532 2089 2540
rect 2066 2528 2070 2531
rect 2070 2502 2073 2518
rect 1934 2472 1937 2478
rect 1946 2468 1950 2471
rect 1986 2468 1990 2471
rect 2018 2468 2022 2471
rect 1974 2462 1977 2468
rect 2054 2462 2057 2498
rect 2078 2492 2081 2508
rect 2102 2492 2105 2518
rect 2070 2482 2073 2488
rect 2078 2482 2081 2488
rect 2106 2478 2110 2481
rect 2134 2481 2137 2658
rect 2182 2652 2185 2658
rect 2222 2642 2225 2658
rect 2230 2612 2233 2668
rect 2310 2661 2313 2918
rect 2318 2842 2321 2898
rect 2374 2892 2377 2918
rect 2446 2912 2449 3038
rect 2454 2952 2457 3048
rect 2510 3042 2513 3078
rect 2518 3052 2521 3058
rect 2526 3041 2529 3068
rect 2550 3061 2553 3118
rect 2582 3112 2585 3138
rect 2582 3072 2585 3108
rect 2590 3092 2593 3218
rect 2638 3192 2641 3248
rect 2654 3242 2657 3268
rect 2666 3258 2670 3261
rect 2698 3258 2702 3261
rect 2710 3231 2713 3258
rect 2766 3251 2769 3328
rect 2798 3292 2801 3328
rect 2814 3302 2817 3328
rect 2926 3302 2929 3328
rect 2814 3272 2817 3278
rect 2774 3262 2777 3268
rect 2766 3248 2777 3251
rect 2722 3238 2726 3241
rect 2710 3228 2721 3231
rect 2718 3192 2721 3228
rect 2774 3192 2777 3248
rect 2782 3232 2785 3268
rect 2854 3262 2857 3268
rect 2826 3258 2830 3261
rect 2842 3258 2846 3261
rect 2670 3172 2673 3178
rect 2702 3162 2705 3168
rect 2710 3162 2713 3168
rect 2646 3152 2649 3158
rect 2678 3142 2681 3158
rect 2798 3152 2801 3258
rect 2886 3252 2889 3259
rect 2822 3248 2830 3251
rect 2850 3248 2854 3251
rect 2822 3222 2825 3248
rect 2830 3152 2833 3238
rect 2894 3232 2897 3268
rect 2894 3152 2897 3228
rect 2934 3192 2937 3298
rect 2942 3262 2945 3328
rect 2958 3302 2961 3328
rect 2974 3292 2977 3328
rect 2998 3292 3001 3328
rect 3022 3292 3025 3328
rect 3062 3328 3066 3332
rect 3086 3328 3090 3332
rect 3110 3331 3114 3332
rect 3158 3331 3162 3332
rect 3102 3328 3114 3331
rect 3150 3328 3162 3331
rect 3182 3331 3186 3332
rect 3206 3331 3210 3332
rect 3230 3331 3234 3332
rect 3326 3331 3330 3332
rect 3350 3331 3354 3332
rect 3182 3328 3193 3331
rect 3206 3328 3217 3331
rect 3230 3328 3241 3331
rect 3040 3303 3042 3307
rect 3046 3303 3049 3307
rect 3053 3303 3056 3307
rect 3062 3292 3065 3328
rect 3086 3302 3089 3328
rect 2950 3282 2953 3288
rect 2982 3262 2985 3278
rect 2654 3132 2657 3138
rect 2686 3132 2689 3148
rect 2734 3142 2737 3148
rect 2750 3132 2753 3148
rect 2782 3142 2785 3148
rect 2890 3148 2894 3151
rect 2790 3132 2793 3138
rect 2810 3128 2814 3131
rect 2562 3068 2566 3071
rect 2654 3062 2657 3068
rect 2550 3058 2561 3061
rect 2518 3038 2529 3041
rect 2518 3032 2521 3038
rect 2526 2992 2529 3028
rect 2536 3003 2538 3007
rect 2542 3003 2545 3007
rect 2549 3003 2552 3007
rect 2558 2972 2561 3058
rect 2646 3058 2654 3061
rect 2574 3022 2577 3058
rect 2582 3048 2590 3051
rect 2462 2962 2465 2968
rect 2558 2962 2561 2968
rect 2518 2952 2521 2958
rect 2542 2952 2545 2958
rect 2582 2952 2585 3048
rect 2458 2928 2462 2931
rect 2478 2922 2481 2948
rect 2390 2882 2393 2888
rect 2398 2882 2401 2888
rect 2446 2882 2449 2908
rect 2486 2892 2489 2938
rect 2494 2932 2497 2948
rect 2514 2938 2518 2941
rect 2526 2931 2529 2948
rect 2518 2928 2529 2931
rect 2606 2932 2609 2948
rect 2502 2902 2505 2918
rect 2518 2892 2521 2928
rect 2622 2892 2625 3058
rect 2630 3052 2633 3058
rect 2646 2942 2649 3058
rect 2670 3042 2673 3128
rect 2702 3122 2705 3128
rect 2750 3112 2753 3128
rect 2686 3092 2689 3108
rect 2798 3092 2801 3128
rect 2862 3122 2865 3147
rect 2838 3092 2841 3118
rect 2858 3078 2862 3081
rect 2702 3072 2705 3078
rect 2718 3052 2721 3059
rect 2686 2952 2689 3018
rect 2710 2952 2713 2998
rect 2718 2992 2721 3038
rect 2750 2992 2753 3058
rect 2782 3022 2785 3068
rect 2810 3058 2814 3061
rect 2822 3052 2825 3058
rect 2830 3022 2833 3068
rect 2870 3062 2873 3118
rect 2886 3072 2889 3148
rect 2926 3122 2929 3168
rect 2958 3162 2961 3258
rect 3006 3252 3009 3258
rect 3030 3242 3033 3258
rect 2970 3178 2974 3181
rect 3054 3162 3057 3248
rect 3070 3242 3073 3278
rect 3086 3252 3089 3258
rect 3094 3252 3097 3258
rect 3082 3238 3086 3241
rect 2974 3152 2977 3158
rect 2958 3132 2961 3148
rect 2922 3118 2926 3121
rect 2914 3058 2918 3061
rect 2734 2952 2737 2978
rect 2662 2932 2665 2948
rect 2734 2942 2737 2948
rect 2666 2928 2670 2931
rect 2690 2928 2694 2931
rect 2722 2918 2726 2921
rect 2430 2872 2433 2878
rect 2378 2868 2382 2871
rect 2450 2868 2454 2871
rect 2326 2852 2329 2858
rect 2334 2852 2337 2858
rect 2326 2822 2329 2828
rect 2358 2752 2361 2858
rect 2366 2802 2369 2848
rect 2406 2842 2409 2868
rect 2414 2862 2417 2868
rect 2422 2862 2425 2868
rect 2462 2862 2465 2888
rect 2502 2872 2505 2888
rect 2526 2872 2529 2878
rect 2534 2872 2537 2888
rect 2630 2882 2633 2888
rect 2594 2878 2598 2881
rect 2638 2872 2641 2878
rect 2646 2872 2649 2898
rect 2670 2872 2673 2918
rect 2694 2892 2697 2918
rect 2750 2892 2753 2918
rect 2758 2892 2761 3018
rect 2782 3002 2785 3018
rect 2798 2932 2801 3018
rect 2806 2942 2809 3008
rect 2846 2992 2849 3058
rect 2950 2992 2953 3058
rect 2934 2962 2937 2968
rect 2834 2958 2838 2961
rect 2870 2952 2873 2958
rect 2898 2948 2902 2951
rect 2946 2948 2950 2951
rect 2814 2912 2817 2938
rect 2774 2892 2777 2908
rect 2822 2902 2825 2918
rect 2726 2872 2729 2878
rect 2474 2868 2478 2871
rect 2490 2868 2494 2871
rect 2570 2868 2574 2871
rect 2706 2868 2710 2871
rect 2498 2858 2502 2861
rect 2554 2858 2558 2861
rect 2602 2858 2606 2861
rect 2366 2792 2369 2798
rect 2422 2782 2425 2858
rect 2582 2852 2585 2858
rect 2450 2848 2454 2851
rect 2474 2848 2478 2851
rect 2438 2792 2441 2828
rect 2574 2812 2577 2848
rect 2614 2832 2617 2868
rect 2638 2862 2641 2868
rect 2686 2862 2689 2868
rect 2702 2852 2705 2858
rect 2662 2842 2665 2848
rect 2674 2838 2678 2841
rect 2686 2832 2689 2848
rect 2694 2822 2697 2848
rect 2486 2792 2489 2808
rect 2536 2803 2538 2807
rect 2542 2803 2545 2807
rect 2549 2803 2552 2807
rect 2342 2742 2345 2748
rect 2334 2732 2337 2738
rect 2350 2732 2353 2738
rect 2326 2721 2329 2728
rect 2326 2718 2337 2721
rect 2318 2681 2321 2718
rect 2318 2678 2329 2681
rect 2318 2662 2321 2668
rect 2306 2658 2318 2661
rect 2326 2652 2329 2678
rect 2262 2582 2265 2618
rect 2150 2542 2153 2568
rect 2166 2542 2169 2558
rect 2174 2542 2177 2568
rect 2194 2558 2201 2561
rect 2190 2542 2193 2548
rect 2158 2532 2161 2538
rect 2186 2528 2190 2531
rect 2198 2522 2201 2558
rect 2262 2552 2265 2558
rect 2286 2552 2289 2558
rect 2218 2548 2222 2551
rect 2282 2548 2286 2551
rect 2294 2542 2297 2548
rect 2242 2538 2249 2541
rect 2210 2528 2214 2531
rect 2158 2492 2161 2508
rect 2174 2492 2177 2518
rect 2126 2478 2137 2481
rect 2206 2482 2209 2488
rect 2086 2472 2089 2478
rect 2126 2472 2129 2478
rect 2066 2468 2070 2471
rect 1958 2422 1961 2448
rect 2086 2442 2089 2468
rect 2230 2462 2233 2468
rect 2134 2452 2137 2458
rect 2190 2452 2193 2458
rect 2222 2452 2225 2458
rect 2102 2442 2105 2448
rect 2158 2442 2161 2448
rect 1886 2392 1889 2408
rect 1926 2392 1929 2418
rect 2070 2392 2073 2408
rect 2094 2372 2097 2418
rect 2066 2368 2070 2371
rect 1746 2358 1750 2361
rect 1718 2342 1721 2358
rect 1734 2342 1737 2348
rect 1766 2342 1769 2348
rect 1774 2342 1777 2368
rect 1846 2358 1865 2361
rect 1798 2352 1801 2358
rect 1782 2342 1785 2348
rect 1822 2342 1825 2348
rect 1746 2338 1750 2341
rect 1754 2328 1758 2331
rect 1778 2328 1782 2331
rect 1718 2272 1721 2278
rect 1726 2272 1729 2298
rect 1742 2272 1745 2278
rect 1750 2272 1753 2298
rect 1706 2268 1713 2271
rect 1698 2248 1702 2251
rect 1662 2172 1665 2248
rect 1670 2162 1673 2178
rect 1654 2152 1657 2158
rect 1618 2148 1622 2151
rect 1578 2138 1582 2141
rect 1634 2138 1638 2141
rect 1678 2141 1681 2218
rect 1710 2212 1713 2268
rect 1746 2248 1750 2251
rect 1766 2251 1769 2298
rect 1782 2272 1785 2278
rect 1766 2248 1774 2251
rect 1790 2251 1793 2308
rect 1798 2292 1801 2338
rect 1846 2332 1849 2358
rect 1842 2328 1846 2331
rect 1854 2331 1857 2348
rect 1862 2342 1865 2358
rect 1854 2328 1862 2331
rect 1866 2328 1870 2331
rect 1830 2312 1833 2328
rect 1814 2282 1817 2288
rect 1802 2278 1806 2281
rect 1830 2272 1833 2298
rect 1842 2288 1846 2291
rect 1842 2278 1846 2281
rect 1878 2272 1881 2278
rect 1822 2252 1825 2258
rect 1790 2248 1798 2251
rect 1718 2182 1721 2188
rect 1750 2162 1753 2188
rect 1674 2138 1681 2141
rect 1574 2122 1577 2128
rect 1582 2122 1585 2138
rect 1566 2072 1569 2118
rect 1606 2112 1609 2118
rect 1590 2072 1593 2078
rect 1622 2072 1625 2138
rect 1630 2082 1633 2088
rect 1610 2058 1614 2061
rect 1298 1948 1302 1951
rect 1250 1938 1254 1941
rect 1294 1932 1297 1938
rect 1318 1931 1321 1958
rect 1326 1952 1329 1958
rect 1334 1941 1337 1958
rect 1358 1952 1361 1958
rect 1330 1938 1337 1941
rect 1318 1928 1329 1931
rect 1146 1878 1150 1881
rect 1158 1878 1166 1881
rect 1158 1862 1161 1878
rect 1174 1862 1177 1868
rect 1182 1862 1185 1878
rect 1206 1862 1209 1868
rect 1126 1852 1129 1858
rect 1110 1732 1113 1738
rect 1118 1682 1121 1708
rect 1106 1678 1110 1681
rect 1070 1668 1078 1671
rect 1086 1661 1089 1668
rect 1126 1662 1129 1848
rect 1134 1842 1137 1858
rect 1214 1842 1217 1868
rect 1222 1862 1225 1908
rect 1230 1892 1233 1918
rect 1286 1912 1289 1918
rect 1230 1882 1233 1888
rect 1254 1862 1257 1868
rect 1278 1862 1281 1878
rect 1310 1861 1313 1928
rect 1318 1892 1321 1918
rect 1326 1892 1329 1928
rect 1342 1892 1345 1948
rect 1366 1932 1369 2018
rect 1374 1992 1377 1998
rect 1406 1992 1409 2008
rect 1438 1962 1441 2038
rect 1462 1972 1465 2018
rect 1512 2003 1514 2007
rect 1518 2003 1521 2007
rect 1525 2003 1528 2007
rect 1534 2002 1537 2058
rect 1566 2052 1569 2058
rect 1570 2048 1574 2051
rect 1638 2042 1641 2068
rect 1478 1962 1481 1998
rect 1542 1982 1545 2018
rect 1598 1992 1601 2028
rect 1646 2022 1649 2138
rect 1662 2072 1665 2118
rect 1678 2062 1681 2118
rect 1686 2082 1689 2088
rect 1678 2032 1681 2048
rect 1694 2042 1697 2138
rect 1702 2062 1705 2158
rect 1734 2132 1737 2138
rect 1758 2122 1761 2218
rect 1766 2192 1769 2248
rect 1766 2162 1769 2188
rect 1782 2152 1785 2198
rect 1782 2142 1785 2148
rect 1790 2142 1793 2178
rect 1798 2152 1801 2198
rect 1830 2152 1833 2178
rect 1818 2138 1822 2141
rect 1786 2128 1793 2131
rect 1718 2072 1721 2088
rect 1726 2062 1729 2098
rect 1742 2052 1745 2118
rect 1730 2018 1734 2021
rect 1522 1958 1526 1961
rect 1378 1948 1382 1951
rect 1382 1932 1385 1938
rect 1318 1872 1321 1878
rect 1306 1858 1313 1861
rect 1222 1822 1225 1858
rect 1262 1852 1265 1858
rect 1290 1838 1294 1841
rect 1190 1802 1193 1818
rect 1174 1792 1177 1798
rect 1194 1788 1198 1791
rect 1134 1782 1137 1788
rect 1162 1758 1166 1761
rect 1222 1752 1225 1798
rect 1246 1752 1249 1828
rect 1286 1762 1289 1768
rect 1154 1748 1161 1751
rect 1138 1738 1142 1741
rect 1134 1682 1137 1708
rect 1134 1662 1137 1678
rect 1150 1672 1153 1738
rect 1158 1722 1161 1748
rect 1210 1748 1214 1751
rect 1266 1748 1270 1751
rect 1282 1748 1286 1751
rect 1182 1732 1185 1738
rect 1190 1722 1193 1748
rect 1282 1738 1286 1741
rect 1230 1732 1233 1738
rect 1210 1728 1214 1731
rect 1274 1728 1278 1731
rect 1082 1658 1089 1661
rect 1098 1658 1102 1661
rect 1050 1648 1054 1651
rect 1026 1618 1030 1621
rect 1070 1612 1073 1618
rect 982 1562 985 1568
rect 1006 1542 1009 1608
rect 974 1528 985 1531
rect 958 1508 969 1511
rect 918 1482 921 1508
rect 910 1472 913 1478
rect 942 1472 945 1478
rect 922 1468 926 1471
rect 950 1462 953 1478
rect 942 1458 950 1461
rect 798 1438 809 1441
rect 930 1448 934 1451
rect 726 1361 729 1418
rect 726 1358 734 1361
rect 730 1348 734 1351
rect 742 1342 745 1438
rect 782 1432 785 1438
rect 714 1338 718 1341
rect 742 1322 745 1338
rect 702 1312 705 1318
rect 734 1302 737 1318
rect 750 1302 753 1398
rect 782 1362 785 1368
rect 758 1352 761 1358
rect 790 1352 793 1398
rect 798 1382 801 1438
rect 838 1432 841 1448
rect 874 1438 878 1441
rect 922 1438 926 1441
rect 942 1392 945 1458
rect 810 1388 814 1391
rect 894 1382 897 1388
rect 958 1382 961 1508
rect 974 1491 977 1518
rect 966 1488 977 1491
rect 798 1352 801 1368
rect 702 1292 705 1298
rect 710 1282 713 1298
rect 686 1268 694 1271
rect 722 1268 726 1271
rect 686 1251 689 1258
rect 718 1252 721 1258
rect 686 1248 694 1251
rect 686 1222 689 1228
rect 734 1162 737 1298
rect 742 1272 745 1278
rect 742 1201 745 1218
rect 742 1198 750 1201
rect 638 1102 641 1148
rect 646 1142 649 1148
rect 654 1142 657 1158
rect 690 1148 694 1151
rect 722 1148 726 1151
rect 678 1142 681 1148
rect 742 1142 745 1148
rect 750 1142 753 1148
rect 758 1142 761 1338
rect 774 1232 777 1318
rect 790 1282 793 1348
rect 806 1272 809 1278
rect 822 1272 825 1338
rect 830 1332 833 1348
rect 838 1332 841 1368
rect 846 1282 849 1298
rect 854 1292 857 1368
rect 878 1362 881 1368
rect 862 1342 865 1348
rect 794 1268 798 1271
rect 834 1268 838 1271
rect 782 1262 785 1268
rect 810 1258 814 1261
rect 798 1232 801 1248
rect 782 1212 785 1218
rect 766 1152 769 1158
rect 698 1138 702 1141
rect 650 1058 654 1061
rect 638 1052 641 1058
rect 662 1052 665 1138
rect 686 1132 689 1138
rect 742 1128 750 1131
rect 734 1112 737 1118
rect 670 1062 673 1068
rect 686 1062 689 1078
rect 678 1052 681 1058
rect 622 1028 633 1031
rect 654 1038 662 1041
rect 622 952 625 1028
rect 630 962 633 1018
rect 646 932 649 948
rect 518 872 521 878
rect 378 848 385 851
rect 390 762 393 858
rect 430 852 433 868
rect 406 822 409 848
rect 398 792 401 798
rect 422 792 425 808
rect 446 762 449 858
rect 370 758 374 761
rect 442 758 446 761
rect 258 738 262 741
rect 182 732 185 738
rect 190 721 193 728
rect 182 718 193 721
rect 182 682 185 718
rect 206 702 209 738
rect 230 692 233 728
rect 270 722 273 758
rect 282 748 286 751
rect 294 742 297 758
rect 302 742 305 758
rect 394 748 398 751
rect 254 692 257 698
rect 190 682 193 688
rect 294 672 297 738
rect 122 668 129 671
rect 138 668 142 671
rect 42 548 46 551
rect 46 472 49 548
rect 34 468 38 471
rect 46 462 49 468
rect 38 458 46 461
rect 22 392 25 458
rect 30 412 33 418
rect 6 352 9 358
rect 22 292 25 378
rect 38 352 41 458
rect 54 392 57 588
rect 62 542 65 638
rect 70 552 73 558
rect 62 492 65 518
rect 78 492 81 648
rect 86 592 89 628
rect 102 552 105 558
rect 90 478 94 481
rect 94 462 97 468
rect 86 392 89 448
rect 102 362 105 548
rect 110 492 113 568
rect 126 542 129 668
rect 138 658 142 661
rect 150 632 153 668
rect 178 658 182 661
rect 134 552 137 558
rect 118 392 121 498
rect 134 461 137 548
rect 142 492 145 608
rect 150 592 153 618
rect 166 581 169 648
rect 182 592 185 598
rect 198 592 201 668
rect 214 642 217 658
rect 222 648 230 651
rect 166 578 177 581
rect 130 458 137 461
rect 150 472 153 578
rect 166 552 169 558
rect 150 392 153 468
rect 166 462 169 478
rect 174 472 177 578
rect 214 542 217 548
rect 202 528 206 531
rect 222 492 225 648
rect 230 592 233 628
rect 238 562 241 658
rect 266 648 270 651
rect 254 592 257 648
rect 270 562 273 588
rect 206 472 209 478
rect 230 472 233 518
rect 214 468 222 471
rect 214 461 217 468
rect 210 458 217 461
rect 230 462 233 468
rect 166 452 169 458
rect 182 442 185 448
rect 206 392 209 428
rect 222 412 225 448
rect 246 442 249 538
rect 254 492 257 508
rect 262 482 265 488
rect 270 451 273 518
rect 278 472 281 668
rect 302 662 305 728
rect 318 692 321 748
rect 358 742 361 748
rect 398 738 406 741
rect 318 682 321 688
rect 294 652 297 658
rect 286 642 289 648
rect 286 552 289 558
rect 286 472 289 538
rect 294 522 297 648
rect 302 561 305 658
rect 302 558 310 561
rect 318 542 321 548
rect 326 542 329 738
rect 334 672 337 738
rect 346 718 350 721
rect 358 672 361 738
rect 366 672 369 678
rect 338 658 342 661
rect 374 612 377 738
rect 398 692 401 738
rect 414 732 417 738
rect 390 662 393 678
rect 398 668 406 671
rect 382 642 385 648
rect 390 642 393 648
rect 398 592 401 668
rect 414 662 417 678
rect 414 592 417 618
rect 370 578 374 581
rect 334 572 337 578
rect 422 572 425 758
rect 430 692 433 728
rect 438 672 441 708
rect 454 692 457 838
rect 462 752 465 868
rect 470 802 473 868
rect 510 852 513 858
rect 522 848 526 851
rect 494 842 497 848
rect 480 803 482 807
rect 486 803 489 807
rect 493 803 496 807
rect 502 762 505 778
rect 526 752 529 828
rect 462 742 465 748
rect 466 728 470 731
rect 462 692 465 718
rect 454 652 457 658
rect 462 652 465 658
rect 430 642 433 648
rect 430 592 433 628
rect 342 558 350 561
rect 334 552 337 558
rect 326 531 329 538
rect 318 528 329 531
rect 318 492 321 528
rect 306 478 310 481
rect 326 472 329 488
rect 334 482 337 548
rect 342 492 345 558
rect 358 532 361 538
rect 366 522 369 548
rect 366 472 369 518
rect 382 512 385 558
rect 438 542 441 558
rect 470 552 473 708
rect 478 672 481 748
rect 518 742 521 748
rect 486 682 489 718
rect 498 688 502 691
rect 478 632 481 648
rect 510 642 513 718
rect 534 692 537 878
rect 582 872 585 928
rect 606 922 609 928
rect 630 892 633 918
rect 654 892 657 1038
rect 678 1012 681 1048
rect 694 1022 697 1098
rect 722 1068 726 1071
rect 714 1058 718 1061
rect 706 1018 710 1021
rect 734 1002 737 1108
rect 742 1092 745 1128
rect 758 1072 761 1138
rect 774 1132 777 1188
rect 814 1162 817 1188
rect 794 1158 798 1161
rect 822 1152 825 1268
rect 826 1148 830 1151
rect 806 1142 809 1148
rect 838 1142 841 1258
rect 846 1171 849 1278
rect 862 1271 865 1338
rect 882 1328 886 1331
rect 894 1321 897 1368
rect 966 1362 969 1488
rect 982 1482 985 1528
rect 992 1503 994 1507
rect 998 1503 1001 1507
rect 1005 1503 1008 1507
rect 974 1472 977 1478
rect 1014 1462 1017 1598
rect 1038 1552 1041 1588
rect 1026 1548 1030 1551
rect 1046 1542 1049 1608
rect 1078 1582 1081 1658
rect 1086 1572 1089 1618
rect 1070 1561 1073 1568
rect 1058 1558 1073 1561
rect 1094 1562 1097 1578
rect 1102 1552 1105 1658
rect 1082 1548 1086 1551
rect 1062 1542 1065 1548
rect 1094 1542 1097 1548
rect 1026 1538 1030 1541
rect 1102 1541 1105 1548
rect 1102 1538 1110 1541
rect 1086 1522 1089 1538
rect 1022 1462 1025 1508
rect 1034 1488 1038 1491
rect 974 1432 977 1458
rect 974 1362 977 1388
rect 998 1362 1001 1458
rect 1006 1452 1009 1458
rect 986 1358 990 1361
rect 902 1352 905 1358
rect 926 1352 929 1358
rect 998 1352 1001 1358
rect 1014 1352 1017 1398
rect 914 1338 918 1341
rect 954 1338 958 1341
rect 886 1318 897 1321
rect 878 1312 881 1318
rect 886 1292 889 1318
rect 862 1268 870 1271
rect 874 1258 878 1261
rect 854 1252 857 1258
rect 846 1168 857 1171
rect 846 1152 849 1158
rect 802 1138 806 1141
rect 818 1138 822 1141
rect 786 1128 790 1131
rect 774 1091 777 1118
rect 830 1092 833 1118
rect 766 1088 777 1091
rect 746 1068 750 1071
rect 742 1022 745 1048
rect 670 912 673 928
rect 542 742 545 868
rect 550 852 553 858
rect 566 772 569 858
rect 574 752 577 868
rect 598 862 601 888
rect 626 878 630 881
rect 610 868 614 871
rect 630 862 633 868
rect 622 852 625 858
rect 582 842 585 848
rect 598 832 601 838
rect 614 832 617 838
rect 598 792 601 818
rect 582 772 585 778
rect 570 748 574 751
rect 542 682 545 718
rect 526 672 529 678
rect 550 662 553 748
rect 558 742 561 748
rect 574 742 577 748
rect 566 672 569 738
rect 582 692 585 738
rect 558 662 561 668
rect 518 652 521 658
rect 558 651 561 658
rect 550 648 561 651
rect 534 642 537 648
rect 480 603 482 607
rect 486 603 489 607
rect 493 603 496 607
rect 498 558 502 561
rect 538 558 542 561
rect 418 538 422 541
rect 422 532 425 538
rect 410 528 414 531
rect 390 522 393 528
rect 414 492 417 508
rect 406 472 409 478
rect 354 468 358 471
rect 278 462 281 468
rect 302 462 305 468
rect 390 462 393 468
rect 398 462 401 468
rect 366 452 369 458
rect 266 448 273 451
rect 102 352 105 358
rect 66 348 70 351
rect 170 348 174 351
rect 86 282 89 288
rect 62 262 65 268
rect 134 262 137 348
rect 158 342 161 348
rect 182 342 185 348
rect 194 338 198 341
rect 206 332 209 348
rect 222 341 225 358
rect 230 352 233 418
rect 222 338 233 341
rect 174 292 177 318
rect 166 262 169 268
rect 6 252 9 258
rect 30 252 33 258
rect 70 252 73 258
rect 6 152 9 248
rect 54 172 57 178
rect 70 152 73 248
rect 110 242 113 248
rect 110 182 113 188
rect 134 152 137 258
rect 182 252 185 328
rect 230 292 233 338
rect 210 288 214 291
rect 238 272 241 388
rect 246 332 249 338
rect 254 292 257 448
rect 342 442 345 448
rect 278 392 281 418
rect 310 362 313 438
rect 334 392 337 408
rect 366 392 369 398
rect 382 392 385 458
rect 414 392 417 458
rect 354 358 361 361
rect 262 352 265 358
rect 282 338 286 341
rect 218 268 222 271
rect 230 268 238 271
rect 182 232 185 248
rect 150 192 153 198
rect 182 192 185 218
rect 190 151 193 258
rect 190 148 198 151
rect 6 62 9 148
rect 30 142 33 148
rect 30 62 33 68
rect 38 62 41 148
rect 54 82 57 88
rect 70 62 73 148
rect 134 142 137 148
rect 166 142 169 148
rect 198 142 201 148
rect 98 138 102 141
rect 118 82 121 88
rect 134 62 137 138
rect 214 132 217 138
rect 154 88 158 91
rect 178 79 185 81
rect 174 78 185 79
rect 182 62 185 78
rect 190 62 193 108
rect 42 58 46 61
rect 210 58 214 61
rect 70 52 73 58
rect 102 52 105 58
rect 86 32 89 38
rect 134 -19 137 58
rect 222 52 225 148
rect 230 92 233 268
rect 254 258 262 261
rect 254 251 257 258
rect 250 248 257 251
rect 262 242 265 248
rect 270 222 273 268
rect 294 261 297 298
rect 310 272 313 358
rect 334 342 337 348
rect 346 338 350 341
rect 318 272 321 338
rect 350 292 353 318
rect 358 292 361 358
rect 366 332 369 348
rect 374 332 377 338
rect 366 271 369 328
rect 382 292 385 338
rect 390 322 393 328
rect 398 292 401 358
rect 366 268 374 271
rect 294 258 318 261
rect 278 242 281 258
rect 286 252 289 258
rect 294 172 297 248
rect 318 242 321 248
rect 310 162 313 168
rect 294 158 302 161
rect 246 112 249 118
rect 246 52 249 58
rect 254 51 257 148
rect 282 138 286 141
rect 286 132 289 138
rect 278 102 281 118
rect 270 62 273 98
rect 294 92 297 158
rect 318 152 321 208
rect 310 148 318 151
rect 310 62 313 148
rect 326 92 329 178
rect 334 162 337 258
rect 342 248 350 251
rect 342 131 345 248
rect 358 192 361 268
rect 390 251 393 278
rect 414 272 417 348
rect 410 268 414 271
rect 422 261 425 448
rect 430 432 433 458
rect 438 371 441 538
rect 454 512 457 548
rect 518 542 521 548
rect 454 422 457 508
rect 462 432 465 458
rect 446 382 449 418
rect 470 392 473 518
rect 478 502 481 538
rect 550 522 553 648
rect 558 592 561 608
rect 566 581 569 668
rect 590 662 593 758
rect 614 742 617 818
rect 630 802 633 858
rect 638 762 641 828
rect 622 742 625 748
rect 606 692 609 728
rect 614 672 617 738
rect 622 692 625 698
rect 558 578 569 581
rect 582 632 585 648
rect 582 582 585 628
rect 558 502 561 578
rect 590 562 593 648
rect 606 641 609 658
rect 606 638 614 641
rect 610 618 614 621
rect 622 592 625 648
rect 630 562 633 738
rect 638 662 641 718
rect 646 672 649 748
rect 654 692 657 848
rect 662 832 665 848
rect 678 842 681 938
rect 686 872 689 988
rect 694 962 697 978
rect 698 948 702 951
rect 686 852 689 858
rect 694 852 697 918
rect 702 872 705 878
rect 678 792 681 818
rect 710 751 713 998
rect 750 992 753 1058
rect 766 1052 769 1088
rect 778 1068 782 1071
rect 794 1058 798 1061
rect 758 1022 761 1028
rect 774 992 777 1028
rect 726 942 729 948
rect 734 892 737 958
rect 782 952 785 1058
rect 806 1052 809 1068
rect 814 1052 817 1058
rect 798 1022 801 1048
rect 822 1041 825 1088
rect 846 1072 849 1138
rect 854 1112 857 1168
rect 870 1162 873 1198
rect 878 1142 881 1148
rect 886 1132 889 1158
rect 862 1082 865 1118
rect 878 1092 881 1128
rect 814 1038 825 1041
rect 834 1068 838 1071
rect 886 1071 889 1118
rect 894 1092 897 1278
rect 902 1252 905 1318
rect 926 1272 929 1298
rect 966 1282 969 1318
rect 974 1302 977 1348
rect 1006 1342 1009 1348
rect 986 1338 990 1341
rect 918 1252 921 1258
rect 902 1222 905 1238
rect 934 1202 937 1278
rect 966 1262 969 1268
rect 974 1262 977 1278
rect 982 1272 985 1308
rect 992 1303 994 1307
rect 998 1303 1001 1307
rect 1005 1303 1008 1307
rect 1014 1291 1017 1298
rect 1006 1288 1017 1291
rect 998 1271 1001 1278
rect 990 1268 1001 1271
rect 1006 1272 1009 1288
rect 1022 1282 1025 1428
rect 1030 1422 1033 1478
rect 1054 1472 1057 1518
rect 1062 1462 1065 1518
rect 1070 1462 1073 1478
rect 1102 1462 1105 1538
rect 1118 1502 1121 1538
rect 1126 1522 1129 1618
rect 1134 1562 1137 1568
rect 1142 1532 1145 1668
rect 1150 1622 1153 1628
rect 1138 1518 1142 1521
rect 1134 1492 1137 1498
rect 1150 1462 1153 1598
rect 1158 1552 1161 1698
rect 1166 1652 1169 1718
rect 1174 1662 1177 1668
rect 1214 1662 1217 1668
rect 1222 1662 1225 1668
rect 1230 1662 1233 1698
rect 1294 1692 1297 1798
rect 1302 1762 1305 1858
rect 1334 1832 1337 1848
rect 1342 1842 1345 1848
rect 1350 1772 1353 1918
rect 1358 1872 1361 1908
rect 1390 1892 1393 1958
rect 1470 1952 1473 1958
rect 1542 1952 1545 1958
rect 1410 1948 1414 1951
rect 1554 1948 1558 1951
rect 1422 1942 1425 1948
rect 1414 1892 1417 1938
rect 1438 1931 1441 1938
rect 1430 1928 1441 1931
rect 1446 1932 1449 1938
rect 1462 1932 1465 1938
rect 1430 1912 1433 1928
rect 1426 1878 1430 1881
rect 1370 1868 1374 1871
rect 1366 1812 1369 1858
rect 1358 1762 1361 1768
rect 1366 1762 1369 1808
rect 1346 1758 1353 1761
rect 1350 1752 1353 1758
rect 1306 1748 1310 1751
rect 1330 1738 1334 1741
rect 1322 1728 1326 1731
rect 1266 1668 1270 1671
rect 1202 1658 1206 1661
rect 1274 1658 1278 1661
rect 1174 1552 1177 1598
rect 1158 1462 1161 1528
rect 1166 1512 1169 1538
rect 1174 1532 1177 1538
rect 1174 1481 1177 1518
rect 1190 1492 1193 1618
rect 1198 1531 1201 1658
rect 1222 1602 1225 1658
rect 1254 1622 1257 1658
rect 1290 1648 1294 1651
rect 1238 1592 1241 1608
rect 1246 1602 1249 1618
rect 1262 1611 1265 1618
rect 1254 1608 1265 1611
rect 1254 1591 1257 1608
rect 1246 1588 1257 1591
rect 1278 1591 1281 1648
rect 1302 1601 1305 1718
rect 1326 1682 1329 1698
rect 1358 1681 1361 1758
rect 1374 1752 1377 1858
rect 1390 1842 1393 1878
rect 1438 1871 1441 1918
rect 1438 1868 1446 1871
rect 1426 1858 1430 1861
rect 1398 1812 1401 1858
rect 1438 1832 1441 1858
rect 1462 1852 1465 1858
rect 1450 1818 1454 1821
rect 1386 1778 1390 1781
rect 1366 1742 1369 1748
rect 1390 1741 1393 1758
rect 1422 1752 1425 1818
rect 1446 1792 1449 1808
rect 1442 1758 1446 1761
rect 1402 1748 1406 1751
rect 1414 1742 1417 1748
rect 1390 1738 1398 1741
rect 1382 1692 1385 1738
rect 1358 1678 1369 1681
rect 1326 1672 1329 1678
rect 1342 1672 1345 1678
rect 1318 1662 1321 1668
rect 1358 1662 1361 1668
rect 1366 1662 1369 1678
rect 1374 1672 1377 1678
rect 1390 1672 1393 1678
rect 1398 1662 1401 1738
rect 1406 1672 1409 1708
rect 1422 1682 1425 1728
rect 1430 1692 1433 1738
rect 1454 1722 1457 1768
rect 1462 1752 1465 1808
rect 1470 1771 1473 1948
rect 1494 1942 1497 1948
rect 1542 1942 1545 1948
rect 1554 1938 1558 1941
rect 1570 1938 1574 1941
rect 1478 1882 1481 1918
rect 1502 1912 1505 1938
rect 1534 1931 1537 1938
rect 1534 1928 1542 1931
rect 1554 1928 1558 1931
rect 1490 1888 1494 1891
rect 1550 1882 1553 1888
rect 1490 1868 1494 1871
rect 1518 1862 1521 1868
rect 1530 1858 1534 1861
rect 1486 1792 1489 1858
rect 1502 1842 1505 1858
rect 1494 1838 1502 1841
rect 1470 1768 1481 1771
rect 1470 1741 1473 1758
rect 1462 1738 1473 1741
rect 1478 1742 1481 1768
rect 1486 1742 1489 1748
rect 1438 1692 1441 1708
rect 1462 1692 1465 1738
rect 1414 1672 1417 1678
rect 1334 1652 1337 1658
rect 1322 1648 1326 1651
rect 1350 1632 1353 1658
rect 1294 1598 1305 1601
rect 1334 1601 1337 1618
rect 1334 1598 1345 1601
rect 1278 1588 1289 1591
rect 1206 1552 1209 1568
rect 1222 1562 1225 1568
rect 1230 1552 1233 1588
rect 1246 1552 1249 1588
rect 1206 1542 1209 1548
rect 1198 1528 1209 1531
rect 1198 1512 1201 1518
rect 1174 1478 1185 1481
rect 1182 1472 1185 1478
rect 1138 1458 1142 1461
rect 1170 1458 1174 1461
rect 1030 1362 1033 1418
rect 1062 1382 1065 1458
rect 1094 1452 1097 1458
rect 1062 1352 1065 1358
rect 1042 1338 1046 1341
rect 1054 1332 1057 1348
rect 1038 1292 1041 1318
rect 1014 1272 1017 1278
rect 1038 1272 1041 1278
rect 946 1258 950 1261
rect 974 1231 977 1258
rect 982 1242 985 1258
rect 974 1228 985 1231
rect 958 1201 961 1218
rect 954 1198 961 1201
rect 934 1152 937 1188
rect 910 1142 913 1148
rect 910 1092 913 1118
rect 882 1068 889 1071
rect 814 982 817 1038
rect 802 958 806 961
rect 814 952 817 978
rect 822 952 825 1008
rect 742 948 750 951
rect 810 948 814 951
rect 718 872 721 878
rect 742 872 745 948
rect 758 942 761 948
rect 754 938 758 941
rect 750 872 753 938
rect 782 932 785 938
rect 790 932 793 938
rect 770 868 774 871
rect 722 858 726 861
rect 726 842 729 848
rect 750 842 753 848
rect 774 832 777 848
rect 762 828 766 831
rect 782 802 785 928
rect 830 922 833 1068
rect 838 1062 841 1068
rect 858 1048 862 1051
rect 850 948 854 951
rect 858 938 862 941
rect 870 932 873 1018
rect 878 962 881 1048
rect 886 1032 889 1058
rect 918 1052 921 1138
rect 942 1132 945 1148
rect 950 1142 953 1188
rect 966 1152 969 1158
rect 970 1138 974 1141
rect 926 1122 929 1128
rect 926 1062 929 1098
rect 942 1072 945 1118
rect 950 1112 953 1138
rect 982 1131 985 1228
rect 990 1221 993 1268
rect 1022 1262 1025 1268
rect 990 1218 1001 1221
rect 998 1202 1001 1218
rect 990 1162 993 1188
rect 974 1128 985 1131
rect 1006 1131 1009 1258
rect 1022 1192 1025 1238
rect 1038 1162 1041 1198
rect 1018 1148 1022 1151
rect 1038 1142 1041 1148
rect 1018 1138 1022 1141
rect 1006 1128 1017 1131
rect 974 1122 977 1128
rect 950 1092 953 1108
rect 890 1018 894 1021
rect 902 1012 905 1048
rect 878 942 881 948
rect 878 922 881 938
rect 798 872 801 898
rect 806 892 809 918
rect 806 872 809 878
rect 794 858 798 861
rect 814 852 817 858
rect 822 851 825 888
rect 830 882 833 918
rect 838 892 841 918
rect 882 888 886 891
rect 834 858 838 861
rect 850 858 854 861
rect 874 858 878 861
rect 822 848 830 851
rect 822 832 825 848
rect 846 842 849 858
rect 790 812 793 818
rect 726 792 729 798
rect 806 792 809 808
rect 814 802 817 818
rect 846 792 849 828
rect 742 782 745 788
rect 718 762 721 768
rect 706 748 713 751
rect 742 742 745 748
rect 674 738 678 741
rect 662 732 665 738
rect 694 732 697 738
rect 702 732 705 738
rect 734 732 737 738
rect 718 702 721 728
rect 726 682 729 688
rect 666 668 670 671
rect 646 652 649 668
rect 678 662 681 668
rect 750 662 753 688
rect 758 672 761 768
rect 766 702 769 758
rect 782 752 785 778
rect 814 762 817 768
rect 822 752 825 758
rect 854 752 857 758
rect 862 751 865 818
rect 886 812 889 848
rect 874 768 878 771
rect 886 762 889 798
rect 894 762 897 1008
rect 902 1002 905 1008
rect 910 992 913 1048
rect 926 952 929 1048
rect 934 1022 937 1068
rect 942 1052 945 1068
rect 950 1032 953 1058
rect 942 962 945 998
rect 950 961 953 1018
rect 958 1002 961 1118
rect 966 1052 969 1078
rect 982 1072 985 1118
rect 992 1103 994 1107
rect 998 1103 1001 1107
rect 1005 1103 1008 1107
rect 1014 1092 1017 1128
rect 1022 1092 1025 1108
rect 986 1058 990 1061
rect 974 1022 977 1058
rect 1022 1052 1025 1058
rect 1010 1018 1014 1021
rect 966 1002 969 1018
rect 962 988 966 991
rect 1014 982 1017 998
rect 950 958 969 961
rect 906 948 918 951
rect 954 948 958 951
rect 910 932 913 938
rect 918 892 921 938
rect 926 902 929 948
rect 942 902 945 918
rect 950 912 953 938
rect 966 912 969 958
rect 974 892 977 958
rect 986 948 990 951
rect 986 938 990 941
rect 938 888 942 891
rect 910 872 913 878
rect 902 812 905 858
rect 918 842 921 888
rect 950 862 953 868
rect 926 832 929 858
rect 918 762 921 768
rect 926 762 929 768
rect 902 752 905 758
rect 862 748 886 751
rect 934 751 937 768
rect 950 762 953 838
rect 958 792 961 878
rect 970 858 974 861
rect 966 842 969 848
rect 982 812 985 908
rect 992 903 994 907
rect 998 903 1001 907
rect 1005 903 1008 907
rect 998 871 1001 888
rect 994 868 1001 871
rect 1014 872 1017 978
rect 1030 962 1033 1128
rect 1046 1081 1049 1278
rect 1054 1202 1057 1288
rect 1070 1282 1073 1448
rect 1110 1432 1113 1458
rect 1082 1428 1086 1431
rect 1086 1352 1089 1418
rect 1098 1348 1102 1351
rect 1110 1342 1113 1428
rect 1102 1332 1105 1338
rect 1118 1331 1121 1418
rect 1126 1341 1129 1458
rect 1158 1442 1161 1448
rect 1174 1432 1177 1438
rect 1170 1388 1177 1391
rect 1134 1352 1137 1358
rect 1126 1338 1137 1341
rect 1110 1328 1121 1331
rect 1110 1292 1113 1328
rect 1094 1282 1097 1288
rect 1062 1262 1065 1268
rect 1070 1262 1073 1268
rect 1102 1262 1105 1268
rect 1078 1241 1081 1258
rect 1094 1252 1097 1258
rect 1066 1238 1081 1241
rect 1066 1198 1073 1201
rect 1054 1142 1057 1148
rect 1062 1092 1065 1158
rect 1070 1082 1073 1198
rect 1078 1192 1081 1198
rect 1078 1142 1081 1148
rect 1078 1102 1081 1138
rect 1086 1092 1089 1148
rect 1094 1142 1097 1228
rect 1046 1078 1057 1081
rect 1038 1062 1041 1068
rect 1046 1062 1049 1068
rect 1038 982 1041 1008
rect 1046 1002 1049 1058
rect 1054 992 1057 1078
rect 1086 1072 1089 1078
rect 1102 1062 1105 1178
rect 1118 1131 1121 1318
rect 1126 1302 1129 1328
rect 1134 1312 1137 1338
rect 1150 1332 1153 1338
rect 1158 1292 1161 1358
rect 1174 1342 1177 1388
rect 1182 1352 1185 1468
rect 1190 1422 1193 1468
rect 1198 1452 1201 1458
rect 1182 1332 1185 1348
rect 1190 1332 1193 1368
rect 1206 1352 1209 1528
rect 1218 1488 1222 1491
rect 1218 1468 1222 1471
rect 1230 1462 1233 1538
rect 1254 1532 1257 1558
rect 1262 1552 1265 1588
rect 1262 1532 1265 1538
rect 1278 1532 1281 1578
rect 1286 1562 1289 1588
rect 1294 1532 1297 1598
rect 1302 1571 1305 1588
rect 1318 1572 1321 1588
rect 1302 1568 1313 1571
rect 1310 1561 1313 1568
rect 1310 1558 1329 1561
rect 1326 1552 1329 1558
rect 1342 1561 1345 1598
rect 1342 1558 1353 1561
rect 1334 1552 1337 1558
rect 1318 1542 1321 1548
rect 1306 1538 1310 1541
rect 1282 1528 1286 1531
rect 1274 1478 1278 1481
rect 1262 1471 1265 1478
rect 1286 1472 1289 1518
rect 1302 1492 1305 1518
rect 1302 1472 1305 1478
rect 1310 1472 1313 1528
rect 1262 1468 1278 1471
rect 1226 1458 1230 1461
rect 1314 1458 1318 1461
rect 1246 1452 1249 1458
rect 1254 1422 1257 1458
rect 1278 1448 1286 1451
rect 1278 1442 1281 1448
rect 1238 1362 1241 1378
rect 1214 1358 1222 1361
rect 1214 1352 1217 1358
rect 1226 1348 1233 1351
rect 1242 1348 1246 1351
rect 1230 1341 1233 1348
rect 1230 1338 1241 1341
rect 1214 1332 1217 1338
rect 1198 1322 1201 1328
rect 1166 1282 1169 1318
rect 1154 1278 1161 1281
rect 1158 1272 1161 1278
rect 1130 1268 1134 1271
rect 1126 1192 1129 1258
rect 1142 1252 1145 1258
rect 1126 1152 1129 1168
rect 1150 1161 1153 1268
rect 1174 1262 1177 1268
rect 1158 1182 1161 1258
rect 1170 1248 1174 1251
rect 1170 1228 1177 1231
rect 1158 1172 1161 1178
rect 1150 1158 1161 1161
rect 1146 1148 1150 1151
rect 1110 1128 1121 1131
rect 1110 1082 1113 1128
rect 1118 1112 1121 1118
rect 1118 1072 1121 1088
rect 1114 1068 1118 1071
rect 1126 1062 1129 1068
rect 1098 1058 1102 1061
rect 1062 1052 1065 1058
rect 1070 1052 1073 1058
rect 1134 1051 1137 1148
rect 1158 1092 1161 1158
rect 1166 1132 1169 1218
rect 1174 1182 1177 1228
rect 1182 1192 1185 1258
rect 1190 1232 1193 1298
rect 1222 1292 1225 1328
rect 1206 1282 1209 1288
rect 1218 1278 1222 1281
rect 1214 1242 1217 1258
rect 1222 1232 1225 1268
rect 1210 1218 1214 1221
rect 1230 1221 1233 1248
rect 1222 1218 1233 1221
rect 1198 1181 1201 1218
rect 1190 1178 1201 1181
rect 1190 1162 1193 1178
rect 1206 1162 1209 1168
rect 1174 1152 1177 1158
rect 1198 1148 1206 1151
rect 1182 1142 1185 1148
rect 1142 1082 1145 1088
rect 1174 1072 1177 1078
rect 1174 1062 1177 1068
rect 1190 1062 1193 1128
rect 1126 1048 1137 1051
rect 1154 1048 1158 1051
rect 1034 958 1041 961
rect 1022 912 1025 918
rect 1014 862 1017 868
rect 1030 862 1033 928
rect 1038 892 1041 958
rect 1062 952 1065 968
rect 1046 942 1049 948
rect 1054 932 1057 938
rect 1078 932 1081 978
rect 1086 952 1089 988
rect 1102 962 1105 1008
rect 1110 971 1113 1038
rect 1126 982 1129 1048
rect 1198 1032 1201 1148
rect 1206 1062 1209 1138
rect 1214 1112 1217 1178
rect 1222 1092 1225 1218
rect 1238 1202 1241 1338
rect 1262 1332 1265 1378
rect 1270 1362 1273 1398
rect 1278 1392 1281 1398
rect 1310 1392 1313 1398
rect 1298 1358 1302 1361
rect 1286 1351 1289 1358
rect 1286 1348 1294 1351
rect 1310 1342 1313 1348
rect 1270 1322 1273 1338
rect 1278 1301 1281 1318
rect 1262 1298 1281 1301
rect 1262 1292 1265 1298
rect 1274 1288 1278 1291
rect 1298 1288 1302 1291
rect 1318 1281 1321 1458
rect 1334 1452 1337 1518
rect 1342 1502 1345 1548
rect 1350 1541 1353 1558
rect 1358 1552 1361 1628
rect 1366 1602 1369 1658
rect 1366 1552 1369 1558
rect 1350 1538 1369 1541
rect 1354 1528 1358 1531
rect 1366 1521 1369 1538
rect 1358 1518 1369 1521
rect 1342 1472 1345 1478
rect 1350 1462 1353 1518
rect 1358 1482 1361 1518
rect 1374 1511 1377 1618
rect 1390 1592 1393 1628
rect 1398 1602 1401 1658
rect 1406 1592 1409 1658
rect 1422 1632 1425 1678
rect 1446 1672 1449 1678
rect 1478 1672 1481 1698
rect 1494 1672 1497 1838
rect 1512 1803 1514 1807
rect 1518 1803 1521 1807
rect 1525 1803 1528 1807
rect 1510 1752 1513 1778
rect 1534 1772 1537 1858
rect 1566 1822 1569 1858
rect 1522 1758 1534 1761
rect 1518 1692 1521 1748
rect 1526 1732 1529 1738
rect 1526 1682 1529 1728
rect 1542 1672 1545 1818
rect 1550 1712 1553 1758
rect 1558 1732 1561 1738
rect 1566 1722 1569 1748
rect 1550 1682 1553 1698
rect 1574 1692 1577 1928
rect 1582 1892 1585 1938
rect 1590 1932 1593 1938
rect 1598 1932 1601 1948
rect 1614 1902 1617 2018
rect 1622 1932 1625 1958
rect 1630 1872 1633 1998
rect 1654 1962 1657 2018
rect 1698 2008 1705 2011
rect 1678 1992 1681 2008
rect 1658 1948 1662 1951
rect 1646 1942 1649 1948
rect 1638 1932 1641 1938
rect 1654 1881 1657 1938
rect 1678 1932 1681 1978
rect 1686 1962 1689 1968
rect 1694 1952 1697 1958
rect 1702 1952 1705 2008
rect 1750 1992 1753 2108
rect 1790 2092 1793 2128
rect 1814 2102 1817 2118
rect 1806 2082 1809 2098
rect 1778 2068 1782 2071
rect 1726 1972 1729 1978
rect 1738 1968 1742 1971
rect 1718 1962 1721 1968
rect 1726 1952 1729 1958
rect 1662 1892 1665 1898
rect 1654 1878 1665 1881
rect 1638 1872 1641 1878
rect 1646 1872 1649 1878
rect 1586 1868 1590 1871
rect 1602 1858 1609 1861
rect 1586 1848 1590 1851
rect 1606 1812 1609 1858
rect 1614 1852 1617 1858
rect 1622 1852 1625 1858
rect 1630 1831 1633 1868
rect 1630 1828 1638 1831
rect 1598 1792 1601 1808
rect 1646 1762 1649 1808
rect 1654 1792 1657 1848
rect 1662 1792 1665 1878
rect 1678 1872 1681 1898
rect 1670 1862 1673 1868
rect 1670 1832 1673 1848
rect 1678 1802 1681 1858
rect 1686 1851 1689 1938
rect 1702 1902 1705 1948
rect 1710 1912 1713 1938
rect 1718 1892 1721 1938
rect 1750 1892 1753 1968
rect 1758 1922 1761 2058
rect 1774 2052 1777 2058
rect 1782 2022 1785 2048
rect 1822 2032 1825 2068
rect 1838 2062 1841 2198
rect 1854 2152 1857 2258
rect 1862 2152 1865 2268
rect 1886 2262 1889 2368
rect 1910 2352 1913 2368
rect 1978 2358 1982 2361
rect 1894 2332 1897 2348
rect 1918 2342 1921 2358
rect 1930 2348 1934 2351
rect 1970 2348 1974 2351
rect 2042 2348 2046 2351
rect 1906 2328 1910 2331
rect 1942 2312 1945 2338
rect 1950 2332 1953 2338
rect 1982 2332 1985 2348
rect 1902 2282 1905 2288
rect 1966 2282 1969 2328
rect 1998 2322 2001 2338
rect 2006 2332 2009 2348
rect 2030 2332 2033 2348
rect 2006 2322 2009 2328
rect 1998 2312 2001 2318
rect 1978 2278 1982 2281
rect 1878 2202 1881 2218
rect 1894 2192 1897 2278
rect 1958 2272 1961 2278
rect 1906 2268 1910 2271
rect 1942 2242 1945 2258
rect 1966 2252 1969 2278
rect 1998 2272 2001 2308
rect 2024 2303 2026 2307
rect 2030 2303 2033 2307
rect 2037 2303 2040 2307
rect 2046 2292 2049 2298
rect 2054 2281 2057 2368
rect 2110 2362 2113 2418
rect 2134 2392 2137 2438
rect 2070 2332 2073 2348
rect 2102 2332 2105 2338
rect 2110 2332 2113 2338
rect 2134 2332 2137 2338
rect 2078 2292 2081 2308
rect 2046 2278 2057 2281
rect 2014 2272 2017 2278
rect 2026 2258 2030 2261
rect 1874 2158 1878 2161
rect 1862 2142 1865 2148
rect 1886 2142 1889 2168
rect 1910 2162 1913 2198
rect 1966 2192 1969 2198
rect 1898 2148 1910 2151
rect 1918 2142 1921 2158
rect 1950 2142 1953 2168
rect 1966 2152 1969 2158
rect 1982 2142 1985 2158
rect 1990 2152 1993 2258
rect 2046 2252 2049 2278
rect 2074 2268 2078 2271
rect 2014 2202 2017 2218
rect 2046 2192 2049 2248
rect 2062 2212 2065 2258
rect 2086 2251 2089 2328
rect 2118 2292 2121 2328
rect 2142 2322 2145 2358
rect 2150 2292 2153 2398
rect 2158 2362 2161 2368
rect 2182 2342 2185 2438
rect 2190 2362 2193 2448
rect 2230 2441 2233 2458
rect 2222 2438 2233 2441
rect 2238 2452 2241 2468
rect 2238 2442 2241 2448
rect 2198 2362 2201 2388
rect 2158 2292 2161 2338
rect 2166 2332 2169 2338
rect 2182 2312 2185 2338
rect 2198 2292 2201 2348
rect 2214 2342 2217 2408
rect 2222 2352 2225 2438
rect 2246 2422 2249 2538
rect 2258 2528 2262 2531
rect 2254 2482 2257 2498
rect 2258 2468 2262 2471
rect 2270 2452 2273 2458
rect 2258 2438 2262 2441
rect 2278 2372 2281 2518
rect 2286 2492 2289 2518
rect 2302 2492 2305 2608
rect 2310 2572 2313 2618
rect 2310 2472 2313 2538
rect 2326 2532 2329 2578
rect 2334 2562 2337 2718
rect 2358 2702 2361 2748
rect 2374 2742 2377 2778
rect 2414 2752 2417 2758
rect 2382 2742 2385 2748
rect 2430 2742 2433 2778
rect 2446 2762 2449 2788
rect 2566 2782 2569 2788
rect 2502 2762 2505 2768
rect 2466 2758 2470 2761
rect 2554 2758 2558 2761
rect 2438 2722 2441 2728
rect 2430 2692 2433 2708
rect 2446 2692 2449 2758
rect 2478 2748 2486 2751
rect 2514 2748 2518 2751
rect 2454 2742 2457 2748
rect 2462 2742 2465 2748
rect 2478 2692 2481 2748
rect 2526 2742 2529 2758
rect 2498 2738 2502 2741
rect 2382 2682 2385 2688
rect 2398 2682 2401 2688
rect 2354 2678 2358 2681
rect 2502 2681 2505 2718
rect 2498 2678 2505 2681
rect 2550 2702 2553 2748
rect 2550 2682 2553 2698
rect 2342 2662 2345 2668
rect 2346 2618 2350 2621
rect 2366 2592 2369 2678
rect 2402 2668 2406 2671
rect 2418 2666 2422 2669
rect 2382 2592 2385 2638
rect 2342 2542 2345 2558
rect 2350 2552 2353 2558
rect 2406 2552 2409 2598
rect 2430 2592 2433 2618
rect 2438 2572 2441 2678
rect 2494 2672 2497 2678
rect 2462 2662 2465 2668
rect 2470 2652 2473 2668
rect 2502 2661 2505 2668
rect 2534 2662 2537 2668
rect 2498 2658 2505 2661
rect 2514 2658 2518 2661
rect 2470 2642 2473 2648
rect 2526 2642 2529 2658
rect 2498 2558 2502 2561
rect 2354 2538 2358 2541
rect 2326 2492 2329 2528
rect 2374 2512 2377 2528
rect 2390 2512 2393 2528
rect 2398 2522 2401 2528
rect 2398 2492 2401 2508
rect 2342 2482 2345 2488
rect 2406 2482 2409 2528
rect 2414 2492 2417 2558
rect 2438 2542 2441 2548
rect 2438 2522 2441 2538
rect 2346 2468 2350 2471
rect 2434 2468 2438 2471
rect 2318 2462 2321 2468
rect 2286 2442 2289 2448
rect 2294 2442 2297 2448
rect 2318 2412 2321 2458
rect 2326 2452 2329 2468
rect 2358 2452 2361 2458
rect 2366 2452 2369 2458
rect 2326 2392 2329 2448
rect 2374 2442 2377 2448
rect 2346 2438 2350 2441
rect 2374 2392 2377 2408
rect 2382 2402 2385 2458
rect 2390 2412 2393 2468
rect 2406 2392 2409 2468
rect 2446 2462 2449 2558
rect 2454 2492 2457 2558
rect 2486 2552 2489 2558
rect 2518 2552 2521 2618
rect 2526 2602 2529 2638
rect 2536 2603 2538 2607
rect 2542 2603 2545 2607
rect 2549 2603 2552 2607
rect 2558 2572 2561 2668
rect 2566 2662 2569 2748
rect 2574 2672 2577 2738
rect 2582 2682 2585 2748
rect 2578 2658 2582 2661
rect 2578 2638 2582 2641
rect 2590 2611 2593 2818
rect 2598 2732 2601 2768
rect 2686 2762 2689 2778
rect 2670 2752 2673 2758
rect 2598 2712 2601 2728
rect 2614 2722 2617 2728
rect 2630 2722 2633 2748
rect 2638 2742 2641 2748
rect 2654 2732 2657 2748
rect 2662 2742 2665 2748
rect 2598 2672 2601 2698
rect 2606 2662 2609 2678
rect 2614 2662 2617 2698
rect 2646 2692 2649 2698
rect 2634 2688 2638 2691
rect 2654 2682 2657 2698
rect 2638 2672 2641 2678
rect 2662 2672 2665 2708
rect 2670 2692 2673 2718
rect 2622 2662 2625 2668
rect 2590 2608 2598 2611
rect 2606 2592 2609 2658
rect 2586 2578 2590 2581
rect 2614 2572 2617 2578
rect 2474 2538 2478 2541
rect 2490 2538 2494 2541
rect 2462 2502 2465 2538
rect 2482 2518 2486 2521
rect 2510 2512 2513 2548
rect 2526 2532 2529 2538
rect 2454 2482 2457 2488
rect 2454 2472 2457 2478
rect 2414 2432 2417 2448
rect 2438 2432 2441 2458
rect 2234 2368 2238 2371
rect 2342 2368 2366 2371
rect 2270 2361 2273 2368
rect 2286 2361 2289 2368
rect 2270 2358 2289 2361
rect 2234 2348 2241 2351
rect 2198 2282 2201 2288
rect 2126 2272 2129 2278
rect 2142 2272 2145 2278
rect 2106 2268 2110 2271
rect 2134 2262 2137 2268
rect 2082 2248 2089 2251
rect 2110 2212 2113 2248
rect 2006 2142 2009 2158
rect 2030 2152 2033 2168
rect 1850 2138 1854 2141
rect 1962 2138 1966 2141
rect 1970 2138 1977 2141
rect 1918 2132 1921 2138
rect 1974 2131 1977 2138
rect 1990 2131 1993 2138
rect 1974 2128 1993 2131
rect 1846 2062 1849 2118
rect 1862 2092 1865 2098
rect 1782 1962 1785 1998
rect 1766 1932 1769 1938
rect 1774 1922 1777 1928
rect 1782 1922 1785 1928
rect 1782 1892 1785 1908
rect 1790 1881 1793 1998
rect 1830 1982 1833 2058
rect 1854 2042 1857 2078
rect 1870 2051 1873 2118
rect 1878 2082 1881 2118
rect 1886 2071 1889 2098
rect 1926 2092 1929 2098
rect 1922 2078 1926 2081
rect 1942 2072 1945 2118
rect 1958 2092 1961 2108
rect 1974 2082 1977 2118
rect 2006 2072 2009 2118
rect 2014 2092 2017 2118
rect 2024 2103 2026 2107
rect 2030 2103 2033 2107
rect 2037 2103 2040 2107
rect 1882 2068 1889 2071
rect 2018 2068 2022 2071
rect 1890 2058 1894 2061
rect 1910 2052 1913 2058
rect 1870 2048 1878 2051
rect 1862 2042 1865 2048
rect 1902 2042 1905 2048
rect 1846 1982 1849 2018
rect 1870 1992 1873 2008
rect 1910 1992 1913 2018
rect 1934 2012 1937 2068
rect 1942 2052 1945 2058
rect 1950 2022 1953 2068
rect 1966 2022 1969 2048
rect 1982 2042 1985 2068
rect 1998 2051 2001 2068
rect 1998 2048 2006 2051
rect 1950 1992 1953 1998
rect 1862 1962 1865 1968
rect 1878 1962 1881 1978
rect 1958 1972 1961 1978
rect 1842 1958 1846 1961
rect 1938 1958 1942 1961
rect 1950 1952 1953 1958
rect 1850 1948 1854 1951
rect 1938 1948 1942 1951
rect 1798 1932 1801 1948
rect 1818 1938 1825 1941
rect 1822 1932 1825 1938
rect 1838 1941 1841 1948
rect 1862 1941 1865 1948
rect 1838 1938 1865 1941
rect 1798 1902 1801 1928
rect 1814 1922 1817 1928
rect 1822 1912 1825 1918
rect 1830 1902 1833 1938
rect 1894 1932 1897 1948
rect 1966 1942 1969 2008
rect 1998 1961 2001 2018
rect 2038 1992 2041 2038
rect 1998 1958 2009 1961
rect 1994 1948 1998 1951
rect 1902 1932 1905 1938
rect 1926 1932 1929 1938
rect 1974 1932 1977 1938
rect 1878 1922 1881 1928
rect 1910 1922 1913 1928
rect 1782 1878 1793 1881
rect 1710 1862 1713 1868
rect 1750 1862 1753 1868
rect 1698 1858 1702 1861
rect 1730 1858 1734 1861
rect 1686 1848 1697 1851
rect 1706 1848 1710 1851
rect 1654 1762 1657 1768
rect 1586 1758 1590 1761
rect 1618 1758 1622 1761
rect 1638 1752 1641 1758
rect 1678 1752 1681 1798
rect 1626 1748 1630 1751
rect 1582 1742 1585 1748
rect 1590 1742 1593 1748
rect 1598 1732 1601 1748
rect 1606 1692 1609 1738
rect 1630 1702 1633 1738
rect 1638 1732 1641 1738
rect 1430 1662 1433 1668
rect 1470 1662 1473 1668
rect 1550 1662 1553 1678
rect 1566 1662 1569 1668
rect 1454 1632 1457 1648
rect 1430 1592 1433 1598
rect 1402 1558 1406 1561
rect 1414 1552 1417 1588
rect 1366 1508 1377 1511
rect 1366 1492 1369 1508
rect 1382 1462 1385 1538
rect 1390 1492 1393 1538
rect 1398 1532 1401 1548
rect 1422 1542 1425 1558
rect 1410 1538 1414 1541
rect 1342 1421 1345 1458
rect 1366 1452 1369 1458
rect 1374 1451 1377 1458
rect 1390 1451 1393 1488
rect 1374 1448 1393 1451
rect 1398 1441 1401 1518
rect 1390 1438 1401 1441
rect 1342 1418 1358 1421
rect 1326 1362 1329 1418
rect 1330 1348 1334 1351
rect 1342 1342 1345 1418
rect 1382 1392 1385 1438
rect 1390 1361 1393 1438
rect 1406 1422 1409 1458
rect 1414 1452 1417 1468
rect 1422 1462 1425 1488
rect 1374 1358 1393 1361
rect 1358 1352 1361 1358
rect 1374 1352 1377 1358
rect 1386 1348 1390 1351
rect 1350 1342 1353 1348
rect 1366 1341 1369 1348
rect 1366 1338 1377 1341
rect 1354 1328 1358 1331
rect 1330 1288 1334 1291
rect 1310 1278 1321 1281
rect 1254 1272 1257 1278
rect 1246 1262 1249 1268
rect 1246 1242 1249 1248
rect 1262 1232 1265 1278
rect 1310 1271 1313 1278
rect 1350 1272 1353 1318
rect 1302 1268 1313 1271
rect 1286 1262 1289 1268
rect 1282 1258 1286 1261
rect 1262 1192 1265 1228
rect 1278 1192 1281 1248
rect 1294 1242 1297 1258
rect 1302 1231 1305 1268
rect 1310 1252 1313 1258
rect 1286 1228 1305 1231
rect 1238 1152 1241 1178
rect 1286 1162 1289 1228
rect 1298 1218 1305 1221
rect 1302 1191 1305 1218
rect 1310 1202 1313 1218
rect 1318 1202 1321 1268
rect 1326 1222 1329 1248
rect 1334 1242 1337 1268
rect 1342 1262 1345 1268
rect 1350 1252 1353 1260
rect 1302 1188 1310 1191
rect 1250 1158 1254 1161
rect 1230 1142 1233 1148
rect 1234 1128 1238 1131
rect 1246 1082 1249 1148
rect 1226 1068 1233 1071
rect 1242 1068 1246 1071
rect 1262 1071 1265 1158
rect 1278 1132 1281 1148
rect 1286 1142 1289 1148
rect 1294 1142 1297 1148
rect 1302 1142 1305 1148
rect 1286 1102 1289 1138
rect 1326 1122 1329 1188
rect 1334 1141 1337 1218
rect 1342 1152 1345 1248
rect 1358 1222 1361 1328
rect 1374 1292 1377 1338
rect 1382 1292 1385 1328
rect 1390 1272 1393 1298
rect 1350 1182 1353 1188
rect 1366 1172 1369 1258
rect 1390 1232 1393 1258
rect 1390 1202 1393 1208
rect 1390 1162 1393 1198
rect 1398 1152 1401 1418
rect 1414 1361 1417 1418
rect 1406 1358 1417 1361
rect 1406 1342 1409 1358
rect 1422 1351 1425 1458
rect 1430 1452 1433 1458
rect 1438 1381 1441 1628
rect 1446 1562 1449 1568
rect 1462 1552 1465 1558
rect 1446 1392 1449 1548
rect 1454 1532 1457 1538
rect 1470 1481 1473 1588
rect 1478 1572 1481 1628
rect 1486 1582 1489 1658
rect 1534 1652 1537 1658
rect 1558 1652 1561 1658
rect 1518 1632 1521 1648
rect 1512 1603 1514 1607
rect 1518 1603 1521 1607
rect 1525 1603 1528 1607
rect 1478 1562 1481 1568
rect 1494 1552 1497 1598
rect 1522 1558 1526 1561
rect 1478 1542 1481 1548
rect 1486 1532 1489 1538
rect 1502 1532 1505 1558
rect 1522 1538 1526 1541
rect 1478 1492 1481 1518
rect 1494 1481 1497 1508
rect 1470 1478 1481 1481
rect 1454 1462 1457 1468
rect 1470 1462 1473 1468
rect 1478 1452 1481 1478
rect 1486 1478 1497 1481
rect 1486 1472 1489 1478
rect 1498 1468 1502 1471
rect 1466 1448 1470 1451
rect 1486 1442 1489 1458
rect 1518 1452 1521 1518
rect 1534 1492 1537 1628
rect 1582 1612 1585 1678
rect 1598 1672 1601 1688
rect 1614 1662 1617 1678
rect 1558 1552 1561 1558
rect 1566 1542 1569 1578
rect 1578 1558 1582 1561
rect 1578 1548 1582 1551
rect 1542 1532 1545 1538
rect 1550 1522 1553 1528
rect 1538 1478 1561 1481
rect 1558 1472 1561 1478
rect 1546 1468 1550 1471
rect 1566 1471 1569 1508
rect 1574 1492 1577 1508
rect 1582 1481 1585 1518
rect 1590 1492 1593 1658
rect 1598 1592 1601 1658
rect 1618 1648 1622 1651
rect 1630 1582 1633 1698
rect 1638 1682 1641 1728
rect 1646 1722 1649 1728
rect 1670 1722 1673 1738
rect 1678 1732 1681 1738
rect 1678 1692 1681 1728
rect 1662 1682 1665 1688
rect 1638 1662 1641 1678
rect 1686 1672 1689 1808
rect 1694 1731 1697 1848
rect 1710 1762 1713 1778
rect 1718 1771 1721 1858
rect 1766 1852 1769 1868
rect 1730 1778 1734 1781
rect 1718 1768 1737 1771
rect 1702 1732 1705 1758
rect 1726 1742 1729 1748
rect 1694 1728 1702 1731
rect 1702 1701 1705 1718
rect 1734 1711 1737 1768
rect 1742 1752 1745 1798
rect 1750 1742 1753 1848
rect 1774 1772 1777 1868
rect 1782 1792 1785 1878
rect 1790 1812 1793 1848
rect 1798 1802 1801 1858
rect 1770 1758 1774 1761
rect 1742 1722 1745 1738
rect 1750 1712 1753 1728
rect 1774 1722 1777 1738
rect 1798 1732 1801 1748
rect 1806 1732 1809 1898
rect 1822 1871 1825 1898
rect 1822 1868 1830 1871
rect 1838 1862 1841 1908
rect 1846 1872 1849 1908
rect 1818 1858 1822 1861
rect 1818 1848 1822 1851
rect 1814 1812 1817 1828
rect 1854 1792 1857 1908
rect 1870 1892 1873 1918
rect 1862 1872 1865 1888
rect 1934 1882 1937 1888
rect 1942 1882 1945 1918
rect 1982 1882 1985 1918
rect 2006 1892 2009 1958
rect 2030 1942 2033 1948
rect 2030 1922 2033 1938
rect 2038 1932 2041 1948
rect 2046 1921 2049 2168
rect 2070 2122 2073 2138
rect 2062 2082 2065 2108
rect 2058 2068 2062 2071
rect 2054 1962 2057 2048
rect 2070 2042 2073 2068
rect 2078 1961 2081 2198
rect 2086 2152 2089 2158
rect 2102 2132 2105 2158
rect 2110 2122 2113 2158
rect 2118 2072 2121 2208
rect 2130 2168 2134 2171
rect 2146 2168 2150 2171
rect 2142 2152 2145 2158
rect 2126 2142 2129 2148
rect 2098 2068 2102 2071
rect 2098 2058 2102 2061
rect 2130 2058 2134 2061
rect 2130 2048 2134 2051
rect 2118 2042 2121 2048
rect 2142 2042 2145 2058
rect 2150 2042 2153 2078
rect 2158 2042 2161 2278
rect 2182 2272 2185 2278
rect 2206 2271 2209 2318
rect 2214 2282 2217 2338
rect 2222 2332 2225 2338
rect 2222 2282 2225 2298
rect 2206 2268 2214 2271
rect 2226 2268 2230 2271
rect 2166 2241 2169 2268
rect 2198 2262 2201 2268
rect 2206 2251 2209 2268
rect 2238 2252 2241 2348
rect 2246 2302 2249 2358
rect 2342 2352 2345 2368
rect 2390 2362 2393 2388
rect 2290 2348 2294 2351
rect 2314 2348 2318 2351
rect 2330 2348 2334 2351
rect 2266 2338 2270 2341
rect 2310 2338 2318 2341
rect 2262 2322 2265 2328
rect 2298 2318 2302 2321
rect 2254 2272 2257 2298
rect 2310 2272 2313 2338
rect 2326 2331 2329 2348
rect 2350 2342 2353 2358
rect 2382 2352 2385 2358
rect 2414 2352 2417 2388
rect 2462 2371 2465 2498
rect 2470 2492 2473 2508
rect 2510 2482 2513 2498
rect 2518 2482 2521 2528
rect 2542 2502 2545 2528
rect 2566 2512 2569 2558
rect 2582 2502 2585 2548
rect 2590 2532 2593 2538
rect 2598 2532 2601 2558
rect 2610 2548 2614 2551
rect 2630 2542 2633 2658
rect 2678 2652 2681 2678
rect 2686 2662 2689 2668
rect 2694 2662 2697 2818
rect 2710 2782 2713 2868
rect 2722 2858 2726 2861
rect 2734 2832 2737 2868
rect 2742 2852 2745 2858
rect 2758 2782 2761 2878
rect 2766 2862 2769 2878
rect 2782 2862 2785 2878
rect 2846 2872 2849 2948
rect 2878 2941 2881 2948
rect 2870 2938 2881 2941
rect 2910 2942 2913 2948
rect 2918 2942 2921 2948
rect 2938 2938 2942 2941
rect 2854 2912 2857 2938
rect 2862 2922 2865 2928
rect 2854 2870 2857 2908
rect 2870 2892 2873 2938
rect 2886 2892 2889 2928
rect 2886 2882 2889 2888
rect 2790 2862 2793 2868
rect 2810 2858 2814 2861
rect 2826 2858 2830 2861
rect 2766 2852 2769 2858
rect 2802 2848 2809 2851
rect 2790 2792 2793 2848
rect 2806 2842 2809 2848
rect 2806 2791 2809 2838
rect 2798 2788 2809 2791
rect 2746 2748 2750 2751
rect 2758 2742 2761 2778
rect 2798 2762 2801 2788
rect 2798 2752 2801 2758
rect 2806 2742 2809 2778
rect 2814 2771 2817 2848
rect 2814 2768 2825 2771
rect 2814 2742 2817 2748
rect 2710 2672 2713 2708
rect 2726 2692 2729 2718
rect 2742 2712 2745 2738
rect 2798 2732 2801 2738
rect 2786 2728 2790 2731
rect 2766 2722 2769 2728
rect 2774 2692 2777 2728
rect 2762 2688 2766 2691
rect 2750 2672 2753 2688
rect 2766 2672 2769 2678
rect 2738 2668 2742 2671
rect 2738 2658 2742 2661
rect 2714 2648 2718 2651
rect 2646 2638 2654 2641
rect 2646 2562 2649 2638
rect 2654 2562 2657 2608
rect 2718 2592 2721 2638
rect 2646 2551 2649 2558
rect 2638 2548 2649 2551
rect 2670 2552 2673 2558
rect 2598 2492 2601 2498
rect 2630 2492 2633 2538
rect 2578 2488 2582 2491
rect 2510 2472 2513 2478
rect 2526 2472 2529 2488
rect 2590 2482 2593 2488
rect 2630 2482 2633 2488
rect 2638 2472 2641 2548
rect 2650 2538 2654 2541
rect 2682 2538 2686 2541
rect 2694 2531 2697 2578
rect 2726 2542 2729 2568
rect 2734 2552 2737 2558
rect 2690 2528 2697 2531
rect 2646 2502 2649 2518
rect 2482 2468 2486 2471
rect 2490 2458 2494 2461
rect 2510 2458 2518 2461
rect 2546 2458 2550 2461
rect 2462 2368 2473 2371
rect 2470 2352 2473 2368
rect 2322 2328 2329 2331
rect 2358 2292 2361 2328
rect 2374 2322 2377 2348
rect 2478 2342 2481 2458
rect 2510 2392 2513 2458
rect 2546 2438 2550 2441
rect 2536 2403 2538 2407
rect 2542 2403 2545 2407
rect 2549 2403 2552 2407
rect 2558 2391 2561 2468
rect 2622 2462 2625 2468
rect 2550 2388 2561 2391
rect 2638 2461 2641 2468
rect 2654 2462 2657 2528
rect 2638 2458 2646 2461
rect 2574 2422 2577 2458
rect 2594 2448 2598 2451
rect 2598 2442 2601 2448
rect 2506 2358 2510 2361
rect 2534 2352 2537 2358
rect 2382 2282 2385 2288
rect 2330 2278 2334 2281
rect 2266 2266 2270 2269
rect 2278 2262 2281 2268
rect 2286 2262 2289 2268
rect 2318 2262 2321 2268
rect 2206 2248 2217 2251
rect 2166 2238 2177 2241
rect 2174 2232 2177 2238
rect 2166 2142 2169 2228
rect 2206 2202 2209 2238
rect 2174 2152 2177 2158
rect 2190 2142 2193 2148
rect 2198 2142 2201 2198
rect 2214 2161 2217 2248
rect 2214 2158 2222 2161
rect 2206 2152 2209 2158
rect 2238 2152 2241 2248
rect 2254 2242 2257 2248
rect 2270 2192 2273 2228
rect 2250 2158 2254 2161
rect 2230 2132 2233 2138
rect 2226 2118 2233 2121
rect 2174 2092 2177 2098
rect 2214 2092 2217 2108
rect 2202 2078 2206 2081
rect 2166 2072 2169 2078
rect 2222 2072 2225 2108
rect 2230 2102 2233 2118
rect 2238 2082 2241 2088
rect 2246 2072 2249 2148
rect 2258 2128 2262 2131
rect 2234 2068 2238 2071
rect 2178 2058 2182 2061
rect 2102 2022 2105 2038
rect 2086 1972 2089 2018
rect 2078 1958 2089 1961
rect 2086 1952 2089 1958
rect 2058 1928 2062 1931
rect 2046 1918 2057 1921
rect 2024 1903 2026 1907
rect 2030 1903 2033 1907
rect 2037 1903 2040 1907
rect 1990 1882 1993 1888
rect 2038 1882 2041 1888
rect 2026 1878 2030 1881
rect 2046 1872 2049 1888
rect 1886 1862 1889 1868
rect 1866 1858 1870 1861
rect 1874 1848 1878 1851
rect 1862 1832 1865 1848
rect 1894 1832 1897 1868
rect 1918 1862 1921 1868
rect 1826 1778 1830 1781
rect 1838 1761 1841 1768
rect 1822 1758 1841 1761
rect 1862 1762 1865 1808
rect 1822 1741 1825 1758
rect 1902 1752 1905 1838
rect 1910 1832 1913 1848
rect 1930 1778 1934 1781
rect 1950 1772 1953 1868
rect 1958 1802 1961 1858
rect 1982 1852 1985 1868
rect 1998 1852 2001 1868
rect 2006 1862 2009 1868
rect 2014 1852 2017 1858
rect 1974 1802 1977 1848
rect 1910 1752 1913 1758
rect 1818 1738 1825 1741
rect 1830 1742 1833 1748
rect 1838 1742 1841 1748
rect 1734 1708 1745 1711
rect 1694 1698 1705 1701
rect 1642 1648 1646 1651
rect 1614 1552 1617 1578
rect 1662 1572 1665 1668
rect 1694 1662 1697 1698
rect 1742 1692 1745 1708
rect 1782 1702 1785 1728
rect 1814 1722 1817 1728
rect 1830 1692 1833 1728
rect 1846 1722 1849 1748
rect 1862 1742 1865 1748
rect 1870 1712 1873 1748
rect 1894 1732 1897 1738
rect 1878 1712 1881 1728
rect 1870 1692 1873 1698
rect 1706 1688 1710 1691
rect 1738 1678 1745 1681
rect 1726 1672 1729 1678
rect 1742 1672 1745 1678
rect 1766 1678 1782 1681
rect 1766 1671 1769 1678
rect 1762 1668 1769 1671
rect 1674 1658 1678 1661
rect 1702 1652 1705 1668
rect 1718 1648 1726 1651
rect 1710 1642 1713 1648
rect 1718 1622 1721 1648
rect 1670 1592 1673 1598
rect 1678 1581 1681 1608
rect 1670 1578 1681 1581
rect 1578 1478 1585 1481
rect 1566 1468 1577 1471
rect 1438 1378 1449 1381
rect 1430 1362 1433 1378
rect 1418 1348 1425 1351
rect 1406 1292 1409 1318
rect 1406 1278 1414 1281
rect 1406 1192 1409 1278
rect 1422 1272 1425 1348
rect 1438 1342 1441 1348
rect 1438 1292 1441 1328
rect 1446 1272 1449 1378
rect 1494 1362 1497 1438
rect 1512 1403 1514 1407
rect 1518 1403 1521 1407
rect 1525 1403 1528 1407
rect 1466 1358 1478 1361
rect 1486 1358 1494 1361
rect 1434 1268 1438 1271
rect 1446 1262 1449 1268
rect 1454 1262 1457 1358
rect 1414 1258 1422 1261
rect 1414 1252 1417 1258
rect 1454 1232 1457 1258
rect 1414 1182 1417 1218
rect 1422 1162 1425 1228
rect 1462 1202 1465 1278
rect 1470 1212 1473 1338
rect 1478 1232 1481 1348
rect 1486 1252 1489 1358
rect 1502 1352 1505 1358
rect 1518 1342 1521 1358
rect 1526 1352 1529 1358
rect 1518 1322 1521 1338
rect 1442 1188 1446 1191
rect 1350 1142 1353 1148
rect 1334 1138 1342 1141
rect 1370 1138 1374 1141
rect 1254 1068 1265 1071
rect 1282 1088 1286 1091
rect 1270 1072 1273 1088
rect 1294 1071 1297 1078
rect 1286 1068 1297 1071
rect 1230 1062 1233 1068
rect 1134 992 1137 1018
rect 1110 968 1121 971
rect 1086 942 1089 948
rect 1110 942 1113 958
rect 1118 952 1121 968
rect 930 748 937 751
rect 982 752 985 798
rect 702 652 705 658
rect 710 648 718 651
rect 726 648 734 651
rect 654 592 657 648
rect 710 642 713 648
rect 594 558 601 561
rect 570 548 574 551
rect 482 488 486 491
rect 506 468 510 471
rect 566 471 569 538
rect 598 492 601 558
rect 606 542 609 548
rect 638 542 641 568
rect 662 552 665 608
rect 678 592 681 638
rect 694 572 697 618
rect 710 592 713 628
rect 714 558 718 561
rect 678 548 686 551
rect 654 542 657 548
rect 614 522 617 538
rect 622 492 625 538
rect 646 522 649 528
rect 638 492 641 498
rect 658 488 662 491
rect 622 472 625 488
rect 562 468 569 471
rect 550 462 553 468
rect 598 462 601 468
rect 538 458 542 461
rect 558 452 561 458
rect 526 442 529 448
rect 518 432 521 438
rect 534 432 537 448
rect 480 403 482 407
rect 486 403 489 407
rect 493 403 496 407
rect 526 392 529 418
rect 558 372 561 438
rect 438 368 449 371
rect 438 322 441 328
rect 446 292 449 368
rect 566 362 569 448
rect 582 432 585 458
rect 598 402 601 448
rect 606 392 609 438
rect 614 412 617 468
rect 634 448 638 451
rect 646 451 649 478
rect 662 472 665 478
rect 642 448 649 451
rect 678 452 681 548
rect 694 492 697 558
rect 702 481 705 528
rect 726 502 729 648
rect 750 572 753 618
rect 766 582 769 668
rect 782 652 785 698
rect 790 582 793 738
rect 798 582 801 738
rect 806 662 809 668
rect 806 572 809 618
rect 814 592 817 728
rect 830 721 833 748
rect 822 718 833 721
rect 822 612 825 718
rect 830 672 833 678
rect 846 672 849 748
rect 890 738 894 741
rect 978 738 982 741
rect 870 732 873 738
rect 942 732 945 738
rect 966 732 969 738
rect 990 731 993 848
rect 998 812 1001 818
rect 1002 758 1006 761
rect 1030 742 1033 858
rect 1038 832 1041 868
rect 1046 842 1049 918
rect 1054 882 1057 888
rect 1070 882 1073 918
rect 1094 892 1097 908
rect 1062 872 1065 878
rect 1102 872 1105 918
rect 1118 872 1121 888
rect 1066 858 1070 861
rect 1114 858 1118 861
rect 1126 861 1129 938
rect 1134 892 1137 958
rect 1154 948 1158 951
rect 1166 892 1169 968
rect 1182 961 1185 1018
rect 1174 958 1185 961
rect 1174 942 1177 958
rect 1190 951 1193 988
rect 1186 948 1193 951
rect 1178 938 1185 941
rect 1158 882 1161 888
rect 1126 858 1137 861
rect 1078 851 1081 858
rect 1094 852 1097 858
rect 1058 848 1081 851
rect 982 728 993 731
rect 870 722 873 728
rect 878 702 881 718
rect 866 678 870 681
rect 838 592 841 668
rect 846 662 849 668
rect 886 662 889 698
rect 918 682 921 688
rect 926 671 929 688
rect 922 668 929 671
rect 894 662 897 668
rect 870 652 873 658
rect 894 632 897 658
rect 918 632 921 658
rect 934 651 937 718
rect 958 712 961 718
rect 958 692 961 698
rect 930 648 937 651
rect 950 642 953 668
rect 962 658 969 661
rect 958 631 961 648
rect 966 642 969 658
rect 974 631 977 708
rect 982 691 985 728
rect 1038 722 1041 738
rect 1002 718 1006 721
rect 992 703 994 707
rect 998 703 1001 707
rect 1005 703 1008 707
rect 1030 692 1033 708
rect 1046 692 1049 828
rect 1070 802 1073 818
rect 1086 792 1089 848
rect 1126 832 1129 848
rect 1118 762 1121 768
rect 1062 752 1065 758
rect 1078 742 1081 758
rect 1126 742 1129 748
rect 1058 738 1062 741
rect 1086 738 1094 741
rect 1070 722 1073 738
rect 982 688 993 691
rect 982 672 985 678
rect 958 628 977 631
rect 882 588 886 591
rect 906 588 910 591
rect 734 562 737 568
rect 766 562 769 568
rect 778 548 782 551
rect 694 478 705 481
rect 686 472 689 478
rect 686 452 689 458
rect 678 392 681 448
rect 694 392 697 478
rect 710 452 713 478
rect 706 448 710 451
rect 546 358 550 361
rect 478 352 481 358
rect 454 332 457 348
rect 494 292 497 358
rect 502 342 505 348
rect 526 342 529 348
rect 546 338 550 341
rect 502 272 505 338
rect 534 312 537 338
rect 566 332 569 358
rect 578 348 582 351
rect 590 342 593 368
rect 634 358 638 361
rect 658 358 662 361
rect 610 348 614 351
rect 698 348 702 351
rect 646 342 649 348
rect 654 342 657 348
rect 534 292 537 298
rect 542 292 545 328
rect 598 312 601 338
rect 574 292 577 308
rect 582 282 585 308
rect 622 292 625 328
rect 466 268 470 271
rect 506 268 510 271
rect 462 262 465 268
rect 422 258 430 261
rect 390 248 398 251
rect 350 158 369 161
rect 350 142 353 158
rect 358 142 361 148
rect 342 128 353 131
rect 350 92 353 128
rect 366 92 369 158
rect 374 122 377 158
rect 342 72 345 88
rect 374 82 377 108
rect 382 72 385 168
rect 390 92 393 118
rect 398 72 401 248
rect 414 142 417 188
rect 414 72 417 138
rect 422 92 425 158
rect 430 152 433 258
rect 454 222 457 258
rect 480 203 482 207
rect 486 203 489 207
rect 493 203 496 207
rect 430 72 433 128
rect 438 122 441 148
rect 446 142 449 198
rect 510 192 513 258
rect 558 252 561 258
rect 530 248 534 251
rect 542 241 545 248
rect 534 238 545 241
rect 534 192 537 238
rect 566 202 569 268
rect 582 212 585 278
rect 618 268 622 271
rect 454 162 457 168
rect 454 112 457 118
rect 462 72 465 178
rect 470 142 473 178
rect 494 92 497 158
rect 510 142 513 148
rect 518 142 521 158
rect 526 142 529 178
rect 546 158 550 161
rect 558 152 561 188
rect 590 182 593 268
rect 622 258 630 261
rect 610 248 614 251
rect 622 242 625 258
rect 630 242 633 248
rect 638 242 641 248
rect 570 168 574 171
rect 598 162 601 218
rect 614 192 617 208
rect 614 152 617 178
rect 630 152 633 168
rect 646 152 649 318
rect 662 272 665 278
rect 670 272 673 288
rect 658 258 662 261
rect 678 261 681 348
rect 710 342 713 408
rect 726 392 729 458
rect 734 442 737 548
rect 742 542 745 548
rect 750 531 753 538
rect 742 528 753 531
rect 742 512 745 528
rect 754 478 758 481
rect 782 472 785 488
rect 762 468 766 471
rect 750 452 753 458
rect 762 448 766 451
rect 750 358 758 361
rect 686 322 689 338
rect 710 332 713 338
rect 742 332 745 348
rect 750 331 753 358
rect 766 352 769 378
rect 774 352 777 448
rect 782 382 785 458
rect 790 392 793 548
rect 838 542 841 558
rect 878 552 881 578
rect 918 562 921 628
rect 946 588 950 591
rect 982 562 985 658
rect 850 548 854 551
rect 798 532 801 538
rect 806 522 809 538
rect 870 532 873 538
rect 806 492 809 508
rect 822 492 825 518
rect 846 492 849 498
rect 866 488 870 491
rect 826 468 830 471
rect 854 462 857 478
rect 878 472 881 548
rect 894 522 897 558
rect 902 542 905 548
rect 882 468 886 471
rect 902 462 905 538
rect 910 472 913 558
rect 926 552 929 558
rect 958 552 961 558
rect 990 552 993 688
rect 1038 682 1041 688
rect 1078 682 1081 688
rect 1086 672 1089 738
rect 1094 732 1097 738
rect 1102 722 1105 738
rect 1134 722 1137 858
rect 1142 772 1145 868
rect 1154 848 1158 851
rect 1150 762 1153 778
rect 1142 732 1145 738
rect 1150 732 1153 748
rect 1006 662 1009 668
rect 1014 632 1017 658
rect 1022 648 1030 651
rect 1022 592 1025 648
rect 1054 642 1057 648
rect 1070 642 1073 668
rect 1086 622 1089 668
rect 1110 652 1113 718
rect 1118 672 1121 678
rect 1126 662 1129 718
rect 1158 692 1161 838
rect 1166 792 1169 878
rect 1182 872 1185 938
rect 1198 932 1201 1018
rect 1206 952 1209 1048
rect 1214 992 1217 1048
rect 1210 948 1214 951
rect 1222 941 1225 1058
rect 1254 1052 1257 1068
rect 1262 1052 1265 1058
rect 1258 1028 1262 1031
rect 1270 992 1273 1068
rect 1278 1031 1281 1048
rect 1286 1042 1289 1068
rect 1302 1061 1305 1098
rect 1318 1092 1321 1118
rect 1294 1058 1305 1061
rect 1326 1061 1329 1118
rect 1334 1072 1337 1078
rect 1342 1072 1345 1138
rect 1414 1132 1417 1138
rect 1422 1132 1425 1158
rect 1438 1142 1441 1148
rect 1350 1128 1358 1131
rect 1350 1092 1353 1128
rect 1366 1102 1369 1128
rect 1398 1092 1401 1098
rect 1374 1072 1377 1088
rect 1382 1062 1385 1068
rect 1326 1058 1350 1061
rect 1294 1052 1297 1058
rect 1278 1028 1289 1031
rect 1262 972 1265 988
rect 1270 952 1273 958
rect 1278 952 1281 1018
rect 1286 952 1289 1028
rect 1310 1022 1313 1058
rect 1318 1012 1321 1048
rect 1314 978 1318 981
rect 1234 948 1238 951
rect 1306 948 1313 951
rect 1214 938 1225 941
rect 1190 882 1193 918
rect 1194 868 1198 871
rect 1182 821 1185 858
rect 1198 832 1201 848
rect 1174 818 1185 821
rect 1174 772 1177 818
rect 1206 812 1209 918
rect 1214 892 1217 938
rect 1226 918 1230 921
rect 1230 872 1233 908
rect 1246 902 1249 948
rect 1254 942 1257 948
rect 1262 942 1265 948
rect 1278 942 1281 948
rect 1286 932 1289 938
rect 1294 932 1297 938
rect 1246 882 1249 888
rect 1270 882 1273 888
rect 1278 871 1281 888
rect 1258 868 1281 871
rect 1166 742 1169 748
rect 1182 742 1185 808
rect 1206 752 1209 758
rect 1214 752 1217 848
rect 1222 832 1225 858
rect 1222 762 1225 788
rect 1238 782 1241 868
rect 1254 842 1257 858
rect 1258 828 1262 831
rect 1246 791 1249 828
rect 1246 788 1257 791
rect 1246 772 1249 778
rect 1230 762 1233 768
rect 1182 712 1185 728
rect 1134 672 1137 688
rect 1142 672 1145 678
rect 1154 658 1161 661
rect 1102 632 1105 638
rect 1042 588 1046 591
rect 1062 562 1065 618
rect 1126 582 1129 658
rect 1150 582 1153 618
rect 1090 558 1094 561
rect 1030 552 1033 558
rect 1070 552 1073 558
rect 1110 552 1113 558
rect 1118 552 1121 558
rect 1142 552 1145 558
rect 1130 548 1134 551
rect 934 541 937 548
rect 926 538 937 541
rect 926 522 929 538
rect 942 531 945 548
rect 934 528 945 531
rect 934 492 937 528
rect 966 512 969 548
rect 1046 542 1049 548
rect 1090 538 1094 541
rect 990 532 993 538
rect 1014 532 1017 538
rect 926 482 929 488
rect 942 482 945 488
rect 874 458 878 461
rect 802 448 806 451
rect 814 372 817 448
rect 838 442 841 458
rect 858 448 862 451
rect 838 392 841 438
rect 846 352 849 358
rect 758 342 761 348
rect 774 342 777 348
rect 750 328 761 331
rect 694 292 697 328
rect 718 322 721 328
rect 726 312 729 328
rect 750 272 753 318
rect 758 292 761 328
rect 774 272 777 328
rect 798 312 801 348
rect 814 332 817 348
rect 782 292 785 308
rect 822 302 825 348
rect 838 292 841 308
rect 854 291 857 378
rect 870 362 873 368
rect 862 312 865 358
rect 878 342 881 368
rect 886 362 889 378
rect 902 372 905 458
rect 918 452 921 478
rect 934 468 942 471
rect 934 392 937 468
rect 958 462 961 478
rect 942 442 945 448
rect 914 358 918 361
rect 934 352 937 358
rect 910 342 913 348
rect 918 342 921 348
rect 890 338 894 341
rect 870 292 873 328
rect 854 288 865 291
rect 850 278 854 281
rect 806 272 809 278
rect 862 272 865 288
rect 910 272 913 338
rect 670 258 681 261
rect 818 268 825 271
rect 898 268 905 271
rect 546 148 550 151
rect 558 112 561 148
rect 482 68 486 71
rect 394 58 433 61
rect 250 48 257 51
rect 262 42 265 48
rect 142 -19 146 -18
rect 134 -22 146 -19
rect 166 -19 169 18
rect 174 -19 178 -18
rect 166 -22 178 -19
rect 198 -19 202 -18
rect 206 -19 209 18
rect 270 12 273 58
rect 310 42 313 58
rect 430 52 433 58
rect 362 48 366 51
rect 438 51 441 68
rect 510 62 513 108
rect 542 72 545 98
rect 574 92 577 138
rect 582 132 585 148
rect 634 138 638 141
rect 658 138 662 141
rect 550 72 553 88
rect 582 72 585 118
rect 622 112 625 138
rect 670 122 673 258
rect 686 251 689 268
rect 694 262 697 268
rect 710 252 713 258
rect 686 248 694 251
rect 718 212 721 268
rect 726 262 729 268
rect 742 262 745 268
rect 726 242 729 248
rect 742 242 745 248
rect 758 242 761 248
rect 678 162 681 198
rect 750 192 753 208
rect 774 182 777 268
rect 798 262 801 268
rect 806 262 809 268
rect 794 258 798 261
rect 762 168 766 171
rect 782 171 785 248
rect 790 192 793 228
rect 774 168 785 171
rect 706 158 710 161
rect 686 142 689 158
rect 726 152 729 158
rect 726 142 729 148
rect 738 138 742 141
rect 622 92 625 98
rect 606 72 609 88
rect 674 68 678 71
rect 542 62 545 68
rect 686 62 689 138
rect 718 132 721 138
rect 766 132 769 138
rect 738 128 742 131
rect 774 92 777 168
rect 806 161 809 248
rect 814 182 817 258
rect 822 212 825 268
rect 902 262 905 268
rect 830 248 838 251
rect 830 192 833 248
rect 846 241 849 248
rect 838 238 849 241
rect 870 242 873 248
rect 838 222 841 238
rect 818 168 825 171
rect 822 162 825 168
rect 806 158 817 161
rect 814 152 817 158
rect 754 88 758 91
rect 718 62 721 88
rect 726 72 729 88
rect 434 48 441 51
rect 482 48 486 51
rect 406 32 409 48
rect 454 32 457 48
rect 442 28 446 31
rect 198 -22 209 -19
rect 286 -18 289 8
rect 480 3 482 7
rect 486 3 489 7
rect 493 3 496 7
rect 286 -22 290 -18
rect 510 -19 513 58
rect 534 12 537 58
rect 558 52 561 58
rect 602 48 606 51
rect 606 -18 609 18
rect 622 12 625 48
rect 638 21 641 58
rect 650 48 654 51
rect 662 22 665 58
rect 670 52 673 58
rect 694 22 697 48
rect 726 42 729 58
rect 766 52 769 68
rect 782 52 785 148
rect 806 142 809 148
rect 790 92 793 108
rect 806 72 809 118
rect 822 112 825 158
rect 838 142 841 178
rect 846 162 849 228
rect 846 131 849 158
rect 838 128 849 131
rect 838 92 841 128
rect 854 92 857 208
rect 886 192 889 238
rect 894 182 897 258
rect 902 232 905 248
rect 866 168 870 171
rect 882 158 886 161
rect 862 152 865 158
rect 862 142 865 148
rect 894 142 897 178
rect 902 162 905 208
rect 918 192 921 318
rect 926 272 929 278
rect 934 272 937 338
rect 942 322 945 338
rect 950 292 953 358
rect 958 292 961 458
rect 966 392 969 508
rect 982 492 985 518
rect 992 503 994 507
rect 998 503 1001 507
rect 1005 503 1008 507
rect 986 478 990 481
rect 978 458 985 461
rect 982 392 985 458
rect 990 452 993 458
rect 1014 452 1017 488
rect 1030 482 1033 538
rect 1094 492 1097 508
rect 1102 492 1105 548
rect 1150 542 1153 548
rect 1050 488 1054 491
rect 1038 472 1041 478
rect 1074 468 1078 471
rect 1062 462 1065 468
rect 1030 452 1033 458
rect 1046 442 1049 448
rect 1002 348 1006 351
rect 966 332 969 348
rect 978 338 982 341
rect 994 328 998 331
rect 992 303 994 307
rect 998 303 1001 307
rect 1005 303 1008 307
rect 1014 272 1017 368
rect 1038 352 1041 358
rect 1046 352 1049 438
rect 1062 392 1065 458
rect 1070 381 1073 458
rect 1086 392 1089 488
rect 1102 472 1105 488
rect 1158 482 1161 658
rect 1166 592 1169 708
rect 1190 662 1193 698
rect 1206 682 1209 738
rect 1246 732 1249 748
rect 1254 742 1257 788
rect 1270 752 1273 758
rect 1278 752 1281 848
rect 1286 762 1289 898
rect 1294 862 1297 908
rect 1302 872 1305 898
rect 1310 862 1313 948
rect 1326 951 1329 1058
rect 1338 1038 1342 1041
rect 1350 1038 1358 1041
rect 1334 962 1337 998
rect 1350 992 1353 1038
rect 1366 1031 1369 1058
rect 1358 1028 1369 1031
rect 1326 948 1337 951
rect 1318 942 1321 948
rect 1318 912 1321 938
rect 1326 872 1329 938
rect 1334 932 1337 948
rect 1350 942 1353 948
rect 1358 942 1361 1028
rect 1382 1022 1385 1058
rect 1390 1022 1393 1068
rect 1366 952 1369 988
rect 1382 942 1385 1018
rect 1406 992 1409 1118
rect 1422 1051 1425 1128
rect 1446 1102 1449 1138
rect 1454 1091 1457 1158
rect 1446 1088 1457 1091
rect 1430 1062 1433 1068
rect 1446 1062 1449 1088
rect 1462 1082 1465 1178
rect 1486 1172 1489 1248
rect 1494 1212 1497 1278
rect 1510 1272 1513 1288
rect 1534 1252 1537 1408
rect 1542 1362 1545 1428
rect 1550 1341 1553 1448
rect 1558 1442 1561 1458
rect 1558 1382 1561 1438
rect 1574 1382 1577 1468
rect 1590 1462 1593 1468
rect 1558 1362 1561 1378
rect 1574 1352 1577 1378
rect 1582 1352 1585 1458
rect 1590 1422 1593 1448
rect 1590 1352 1593 1418
rect 1598 1362 1601 1548
rect 1606 1542 1609 1548
rect 1622 1542 1625 1558
rect 1638 1542 1641 1558
rect 1618 1538 1622 1541
rect 1630 1532 1633 1538
rect 1638 1522 1641 1528
rect 1614 1481 1617 1518
rect 1634 1488 1638 1491
rect 1646 1482 1649 1488
rect 1614 1478 1633 1481
rect 1618 1468 1622 1471
rect 1606 1452 1609 1468
rect 1614 1442 1617 1458
rect 1630 1452 1633 1478
rect 1646 1452 1649 1458
rect 1654 1451 1657 1540
rect 1670 1512 1673 1578
rect 1694 1542 1697 1548
rect 1702 1542 1705 1558
rect 1726 1552 1729 1578
rect 1734 1562 1737 1578
rect 1734 1552 1737 1558
rect 1678 1532 1681 1538
rect 1690 1528 1694 1531
rect 1710 1531 1713 1548
rect 1718 1542 1721 1548
rect 1710 1528 1721 1531
rect 1662 1482 1665 1498
rect 1686 1492 1689 1508
rect 1694 1482 1697 1488
rect 1698 1478 1702 1481
rect 1678 1472 1681 1478
rect 1710 1472 1713 1488
rect 1650 1448 1657 1451
rect 1670 1452 1673 1458
rect 1694 1442 1697 1468
rect 1702 1452 1705 1458
rect 1646 1402 1649 1418
rect 1678 1392 1681 1438
rect 1686 1381 1689 1388
rect 1678 1378 1689 1381
rect 1646 1362 1649 1378
rect 1650 1348 1654 1351
rect 1550 1338 1558 1341
rect 1566 1341 1569 1348
rect 1566 1338 1585 1341
rect 1542 1272 1545 1338
rect 1550 1272 1553 1338
rect 1570 1328 1574 1331
rect 1582 1291 1585 1338
rect 1590 1302 1593 1338
rect 1578 1288 1585 1291
rect 1566 1281 1569 1288
rect 1590 1282 1593 1288
rect 1566 1278 1574 1281
rect 1606 1271 1609 1318
rect 1614 1292 1617 1328
rect 1606 1268 1617 1271
rect 1566 1262 1569 1268
rect 1598 1262 1601 1268
rect 1542 1252 1545 1258
rect 1574 1252 1577 1258
rect 1474 1168 1478 1171
rect 1470 1102 1473 1148
rect 1478 1142 1481 1148
rect 1486 1142 1489 1148
rect 1478 1082 1481 1128
rect 1454 1061 1457 1078
rect 1454 1058 1462 1061
rect 1418 1048 1425 1051
rect 1414 952 1417 968
rect 1430 952 1433 1028
rect 1462 1022 1465 1058
rect 1438 992 1441 998
rect 1446 952 1449 988
rect 1358 922 1361 938
rect 1398 932 1401 948
rect 1418 938 1422 941
rect 1446 932 1449 948
rect 1470 942 1473 948
rect 1386 928 1390 931
rect 1454 922 1457 938
rect 1462 932 1465 938
rect 1478 932 1481 1078
rect 1486 1072 1489 1138
rect 1494 1081 1497 1148
rect 1502 1092 1505 1248
rect 1512 1203 1514 1207
rect 1518 1203 1521 1207
rect 1525 1203 1528 1207
rect 1514 1148 1518 1151
rect 1526 1142 1529 1148
rect 1494 1078 1505 1081
rect 1502 1052 1505 1078
rect 1534 1072 1537 1168
rect 1542 1092 1545 1248
rect 1550 1152 1553 1248
rect 1558 1192 1561 1208
rect 1566 1192 1569 1238
rect 1566 1158 1574 1161
rect 1558 1142 1561 1148
rect 1550 1132 1553 1138
rect 1550 1082 1553 1088
rect 1566 1072 1569 1158
rect 1582 1152 1585 1248
rect 1598 1172 1601 1258
rect 1606 1242 1609 1258
rect 1614 1252 1617 1268
rect 1622 1162 1625 1338
rect 1630 1212 1633 1328
rect 1650 1318 1654 1321
rect 1662 1311 1665 1348
rect 1654 1308 1665 1311
rect 1642 1268 1646 1271
rect 1638 1252 1641 1258
rect 1646 1252 1649 1258
rect 1654 1241 1657 1308
rect 1670 1301 1673 1368
rect 1678 1332 1681 1378
rect 1690 1348 1694 1351
rect 1702 1342 1705 1448
rect 1710 1402 1713 1448
rect 1710 1331 1713 1358
rect 1718 1342 1721 1528
rect 1726 1502 1729 1548
rect 1726 1472 1729 1478
rect 1734 1462 1737 1538
rect 1742 1482 1745 1668
rect 1798 1662 1801 1688
rect 1822 1672 1825 1678
rect 1838 1671 1841 1678
rect 1886 1672 1889 1728
rect 1894 1672 1897 1728
rect 1918 1722 1921 1748
rect 1926 1722 1929 1748
rect 1958 1742 1961 1798
rect 1938 1728 1942 1731
rect 1834 1668 1841 1671
rect 1754 1658 1758 1661
rect 1766 1651 1769 1658
rect 1758 1648 1769 1651
rect 1750 1542 1753 1608
rect 1758 1562 1761 1648
rect 1774 1612 1777 1658
rect 1814 1622 1817 1658
rect 1822 1621 1825 1648
rect 1822 1618 1833 1621
rect 1766 1552 1769 1558
rect 1798 1552 1801 1558
rect 1758 1538 1777 1541
rect 1758 1522 1761 1538
rect 1774 1532 1777 1538
rect 1814 1532 1817 1548
rect 1822 1542 1825 1608
rect 1830 1561 1833 1618
rect 1846 1612 1849 1668
rect 1854 1662 1857 1668
rect 1870 1662 1873 1668
rect 1878 1622 1881 1668
rect 1894 1612 1897 1658
rect 1902 1651 1905 1678
rect 1950 1672 1953 1718
rect 1958 1692 1961 1708
rect 1966 1682 1969 1768
rect 1922 1668 1929 1671
rect 1938 1668 1942 1671
rect 1914 1658 1918 1661
rect 1926 1661 1929 1668
rect 1966 1662 1969 1668
rect 1926 1658 1934 1661
rect 1942 1652 1945 1658
rect 1902 1648 1910 1651
rect 1922 1618 1926 1621
rect 1870 1568 1886 1571
rect 1830 1558 1838 1561
rect 1870 1561 1873 1568
rect 1854 1558 1873 1561
rect 1878 1558 1886 1561
rect 1842 1548 1846 1551
rect 1854 1542 1857 1558
rect 1766 1522 1769 1528
rect 1786 1518 1790 1521
rect 1762 1508 1785 1511
rect 1814 1511 1817 1528
rect 1794 1508 1817 1511
rect 1838 1511 1841 1538
rect 1862 1532 1865 1548
rect 1834 1508 1841 1511
rect 1782 1492 1785 1508
rect 1770 1488 1774 1491
rect 1786 1478 1790 1481
rect 1758 1472 1761 1478
rect 1742 1462 1745 1468
rect 1734 1452 1737 1458
rect 1726 1442 1729 1448
rect 1734 1372 1737 1418
rect 1742 1398 1750 1401
rect 1742 1392 1745 1398
rect 1730 1358 1734 1361
rect 1758 1352 1761 1468
rect 1766 1462 1769 1468
rect 1766 1372 1769 1448
rect 1782 1432 1785 1468
rect 1798 1461 1801 1488
rect 1806 1472 1809 1488
rect 1822 1462 1825 1498
rect 1798 1458 1806 1461
rect 1830 1452 1833 1458
rect 1782 1392 1785 1398
rect 1738 1348 1742 1351
rect 1770 1348 1774 1351
rect 1694 1328 1713 1331
rect 1726 1332 1729 1348
rect 1758 1338 1766 1341
rect 1662 1298 1673 1301
rect 1662 1272 1665 1298
rect 1686 1282 1689 1328
rect 1694 1292 1697 1328
rect 1674 1268 1678 1271
rect 1706 1268 1710 1271
rect 1730 1268 1734 1271
rect 1666 1258 1670 1261
rect 1706 1258 1710 1261
rect 1742 1261 1745 1278
rect 1734 1258 1745 1261
rect 1750 1262 1753 1278
rect 1758 1262 1761 1338
rect 1766 1282 1769 1288
rect 1762 1258 1766 1261
rect 1646 1238 1657 1241
rect 1638 1212 1641 1218
rect 1634 1188 1638 1191
rect 1646 1162 1649 1238
rect 1654 1162 1657 1188
rect 1574 1148 1582 1151
rect 1610 1148 1614 1151
rect 1574 1132 1577 1148
rect 1590 1142 1593 1148
rect 1630 1142 1633 1148
rect 1638 1142 1641 1148
rect 1546 1068 1550 1071
rect 1574 1062 1577 1068
rect 1514 1058 1518 1061
rect 1494 962 1497 1018
rect 1502 1012 1505 1048
rect 1558 1022 1561 1048
rect 1512 1003 1514 1007
rect 1518 1003 1521 1007
rect 1525 1003 1528 1007
rect 1558 1002 1561 1018
rect 1566 992 1569 1028
rect 1514 948 1518 951
rect 1490 918 1494 921
rect 1358 912 1361 918
rect 1366 892 1369 908
rect 1322 858 1326 861
rect 1294 812 1297 818
rect 1302 802 1305 858
rect 1334 852 1337 858
rect 1342 812 1345 868
rect 1350 862 1353 878
rect 1366 852 1369 878
rect 1374 852 1377 918
rect 1398 902 1401 918
rect 1518 912 1521 938
rect 1470 908 1497 911
rect 1406 871 1409 908
rect 1414 892 1417 908
rect 1406 868 1417 871
rect 1386 858 1390 861
rect 1386 848 1390 851
rect 1358 802 1361 838
rect 1398 812 1401 868
rect 1406 852 1409 858
rect 1414 841 1417 868
rect 1422 852 1425 878
rect 1434 868 1438 871
rect 1462 871 1465 908
rect 1458 868 1465 871
rect 1470 872 1473 908
rect 1478 862 1481 888
rect 1486 872 1489 898
rect 1494 882 1497 908
rect 1518 882 1521 908
rect 1534 882 1537 988
rect 1542 952 1545 958
rect 1550 892 1553 948
rect 1574 912 1577 1058
rect 1582 992 1585 1138
rect 1614 1082 1617 1128
rect 1590 1078 1609 1081
rect 1622 1081 1625 1138
rect 1622 1078 1633 1081
rect 1590 1072 1593 1078
rect 1590 1052 1593 1058
rect 1598 992 1601 1068
rect 1606 1062 1609 1078
rect 1630 1072 1633 1078
rect 1606 972 1609 1058
rect 1582 952 1585 968
rect 1614 962 1617 998
rect 1602 948 1606 951
rect 1622 942 1625 1068
rect 1630 1052 1633 1058
rect 1638 1041 1641 1128
rect 1646 1062 1649 1148
rect 1654 1092 1657 1148
rect 1662 1122 1665 1138
rect 1654 1072 1657 1078
rect 1662 1072 1665 1098
rect 1670 1082 1673 1188
rect 1678 1152 1681 1248
rect 1694 1162 1697 1228
rect 1718 1162 1721 1258
rect 1734 1192 1737 1258
rect 1774 1252 1777 1308
rect 1782 1241 1785 1348
rect 1790 1342 1793 1438
rect 1798 1352 1801 1428
rect 1838 1422 1841 1468
rect 1806 1322 1809 1418
rect 1814 1352 1817 1388
rect 1822 1362 1825 1368
rect 1830 1332 1833 1358
rect 1846 1352 1849 1508
rect 1854 1472 1857 1508
rect 1862 1492 1865 1518
rect 1870 1512 1873 1538
rect 1878 1521 1881 1558
rect 1894 1552 1897 1558
rect 1910 1552 1913 1618
rect 1958 1592 1961 1648
rect 1974 1572 1977 1688
rect 1982 1672 1985 1748
rect 1990 1742 1993 1828
rect 2054 1792 2057 1918
rect 2078 1912 2081 1948
rect 2094 1942 2097 1948
rect 2086 1932 2089 1938
rect 2102 1932 2105 2018
rect 2158 1972 2161 2018
rect 2166 1992 2169 2058
rect 2190 2052 2193 2058
rect 2198 1972 2201 2018
rect 2214 1992 2217 2048
rect 2254 2042 2257 2118
rect 2270 2112 2273 2178
rect 2286 2152 2289 2258
rect 2310 2252 2313 2258
rect 2342 2242 2345 2258
rect 2366 2252 2369 2278
rect 2386 2268 2390 2271
rect 2398 2262 2401 2338
rect 2414 2312 2417 2338
rect 2422 2282 2425 2338
rect 2470 2332 2473 2338
rect 2494 2332 2497 2338
rect 2506 2328 2510 2331
rect 2550 2322 2553 2388
rect 2574 2342 2577 2418
rect 2594 2358 2598 2361
rect 2606 2352 2609 2358
rect 2586 2348 2590 2351
rect 2614 2341 2617 2368
rect 2622 2352 2625 2458
rect 2630 2362 2633 2458
rect 2654 2362 2657 2458
rect 2670 2452 2673 2458
rect 2678 2452 2681 2518
rect 2686 2472 2689 2528
rect 2710 2512 2713 2538
rect 2726 2522 2729 2538
rect 2750 2532 2753 2538
rect 2758 2521 2761 2528
rect 2750 2518 2761 2521
rect 2694 2462 2697 2498
rect 2630 2352 2633 2358
rect 2614 2338 2622 2341
rect 2562 2328 2566 2331
rect 2454 2302 2457 2318
rect 2406 2272 2409 2278
rect 2454 2272 2457 2278
rect 2434 2268 2438 2271
rect 2394 2258 2398 2261
rect 2422 2252 2425 2268
rect 2434 2258 2438 2261
rect 2442 2248 2446 2251
rect 2334 2192 2337 2208
rect 2422 2172 2425 2218
rect 2406 2162 2409 2168
rect 2346 2158 2350 2161
rect 2302 2152 2305 2158
rect 2322 2148 2326 2151
rect 2278 2142 2281 2148
rect 2306 2138 2310 2141
rect 2326 2122 2329 2138
rect 2366 2132 2369 2148
rect 2374 2142 2377 2158
rect 2414 2152 2417 2158
rect 2430 2152 2433 2198
rect 2486 2192 2489 2318
rect 2566 2292 2569 2318
rect 2574 2282 2577 2338
rect 2646 2332 2649 2358
rect 2654 2352 2657 2358
rect 2658 2338 2662 2341
rect 2670 2341 2673 2448
rect 2702 2442 2705 2468
rect 2710 2392 2713 2508
rect 2722 2458 2726 2461
rect 2726 2452 2729 2458
rect 2734 2452 2737 2498
rect 2742 2442 2745 2458
rect 2750 2452 2753 2518
rect 2766 2472 2769 2518
rect 2758 2462 2761 2468
rect 2766 2452 2769 2458
rect 2734 2392 2737 2438
rect 2774 2422 2777 2668
rect 2782 2662 2785 2668
rect 2790 2532 2793 2718
rect 2802 2688 2806 2691
rect 2814 2672 2817 2738
rect 2822 2732 2825 2768
rect 2830 2742 2833 2818
rect 2838 2742 2841 2868
rect 2846 2842 2849 2868
rect 2878 2862 2881 2868
rect 2842 2738 2846 2741
rect 2830 2702 2833 2718
rect 2846 2712 2849 2718
rect 2846 2692 2849 2708
rect 2834 2688 2838 2691
rect 2854 2682 2857 2738
rect 2862 2682 2865 2738
rect 2886 2732 2889 2758
rect 2894 2742 2897 2748
rect 2870 2702 2873 2718
rect 2866 2678 2870 2681
rect 2826 2668 2830 2671
rect 2798 2662 2801 2668
rect 2806 2642 2809 2668
rect 2838 2662 2841 2678
rect 2846 2672 2849 2678
rect 2878 2672 2881 2688
rect 2894 2672 2897 2698
rect 2910 2682 2913 2938
rect 2938 2928 2942 2931
rect 2926 2882 2929 2888
rect 2958 2882 2961 3128
rect 2974 3082 2977 3148
rect 3006 3142 3009 3147
rect 2990 3082 2993 3118
rect 3014 3092 3017 3158
rect 3038 3142 3041 3148
rect 3078 3132 3081 3138
rect 3022 3082 3025 3128
rect 3094 3122 3097 3128
rect 3030 3072 3033 3118
rect 3040 3103 3042 3107
rect 3046 3103 3049 3107
rect 3053 3103 3056 3107
rect 2994 3058 2998 3061
rect 3006 3042 3009 3068
rect 3062 3062 3065 3078
rect 3070 3062 3073 3068
rect 3042 3058 3046 3061
rect 3054 3032 3057 3048
rect 2982 3002 2985 3018
rect 2982 2982 2985 2988
rect 2966 2962 2969 2968
rect 3010 2958 3014 2961
rect 2982 2952 2985 2958
rect 2926 2821 2929 2838
rect 2918 2818 2929 2821
rect 2918 2742 2921 2818
rect 2926 2762 2929 2768
rect 2910 2672 2913 2678
rect 2870 2662 2873 2668
rect 2866 2658 2870 2661
rect 2806 2492 2809 2618
rect 2814 2582 2817 2658
rect 2846 2652 2849 2658
rect 2894 2651 2897 2668
rect 2906 2658 2910 2661
rect 2894 2648 2910 2651
rect 2854 2592 2857 2628
rect 2894 2612 2897 2618
rect 2918 2602 2921 2738
rect 2926 2722 2929 2728
rect 2926 2672 2929 2718
rect 2934 2712 2937 2858
rect 2966 2752 2969 2818
rect 2974 2802 2977 2938
rect 3014 2882 3017 2948
rect 3022 2942 3025 2978
rect 3046 2952 3049 2958
rect 3070 2942 3073 3048
rect 3078 2982 3081 3118
rect 3086 3082 3089 3088
rect 3086 2952 3089 2958
rect 3102 2952 3105 3328
rect 3150 3292 3153 3328
rect 3190 3292 3193 3328
rect 3214 3292 3217 3328
rect 3238 3292 3241 3328
rect 3318 3328 3330 3331
rect 3342 3328 3354 3331
rect 3502 3328 3506 3332
rect 3542 3331 3546 3332
rect 3542 3328 3553 3331
rect 3318 3292 3321 3328
rect 3342 3292 3345 3328
rect 3126 3282 3129 3288
rect 3114 3278 3118 3281
rect 3386 3278 3390 3281
rect 3314 3268 3318 3271
rect 3378 3268 3382 3271
rect 3482 3268 3486 3271
rect 3110 3262 3113 3268
rect 3438 3262 3441 3268
rect 3462 3262 3465 3268
rect 3122 3258 3126 3261
rect 3178 3258 3182 3261
rect 3386 3258 3390 3261
rect 3118 3242 3121 3248
rect 3138 3238 3142 3241
rect 3110 3152 3113 3178
rect 3142 3151 3145 3158
rect 3126 3072 3129 3138
rect 3166 3072 3169 3258
rect 3198 3182 3201 3258
rect 3202 3178 3206 3181
rect 3222 3172 3225 3258
rect 3218 3158 3222 3161
rect 3174 3142 3177 3148
rect 3230 3132 3233 3168
rect 3246 3152 3249 3258
rect 3294 3192 3297 3238
rect 3334 3162 3337 3258
rect 3358 3242 3361 3258
rect 3366 3252 3369 3258
rect 3398 3252 3401 3258
rect 3494 3252 3497 3258
rect 3450 3248 3454 3251
rect 3502 3251 3505 3328
rect 3514 3278 3518 3281
rect 3514 3268 3518 3271
rect 3514 3258 3518 3261
rect 3522 3258 3526 3261
rect 3502 3248 3513 3251
rect 3274 3158 3278 3161
rect 3306 3158 3310 3161
rect 3334 3152 3337 3158
rect 3238 3112 3241 3128
rect 3182 3092 3185 3108
rect 3178 3088 3182 3091
rect 3214 3082 3217 3088
rect 3246 3082 3249 3148
rect 3254 3072 3257 3148
rect 3326 3132 3329 3138
rect 3334 3092 3337 3148
rect 3350 3132 3353 3168
rect 3358 3152 3361 3158
rect 3358 3132 3361 3138
rect 3374 3132 3377 3238
rect 3398 3232 3401 3238
rect 3382 3152 3385 3158
rect 3414 3142 3417 3248
rect 3398 3132 3401 3138
rect 3378 3128 3382 3131
rect 3350 3122 3353 3128
rect 3314 3088 3318 3091
rect 3342 3082 3345 3118
rect 3382 3092 3385 3118
rect 3390 3082 3393 3118
rect 3422 3112 3425 3248
rect 3470 3232 3473 3248
rect 3430 3192 3433 3218
rect 3122 3059 3126 3062
rect 3190 3052 3193 3058
rect 3126 2992 3129 3048
rect 3198 3042 3201 3068
rect 3214 3062 3217 3068
rect 3246 3052 3249 3059
rect 3318 3042 3321 3078
rect 3438 3072 3441 3148
rect 3334 3051 3337 3068
rect 3334 3048 3345 3051
rect 3222 2992 3225 3038
rect 3242 2958 3246 2961
rect 3154 2948 3158 2951
rect 3034 2938 3038 2941
rect 3082 2938 3086 2941
rect 3030 2882 3033 2938
rect 3054 2922 3057 2928
rect 3040 2903 3042 2907
rect 3046 2903 3049 2907
rect 3053 2903 3056 2907
rect 3014 2872 3017 2878
rect 3054 2872 3057 2878
rect 2994 2868 2998 2871
rect 3062 2862 3065 2938
rect 3070 2872 3073 2938
rect 3102 2932 3105 2938
rect 3082 2888 3086 2891
rect 3018 2848 3022 2851
rect 2986 2818 2990 2821
rect 3030 2792 3033 2798
rect 2998 2752 3001 2758
rect 3006 2752 3009 2778
rect 3018 2768 3022 2771
rect 2978 2748 2982 2751
rect 3026 2748 3030 2751
rect 2942 2682 2945 2738
rect 2950 2722 2953 2728
rect 2950 2692 2953 2708
rect 2958 2682 2961 2718
rect 2974 2712 2977 2748
rect 2986 2738 2990 2741
rect 2982 2692 2985 2698
rect 2986 2678 2990 2681
rect 2998 2672 3001 2738
rect 3010 2668 3014 2671
rect 2814 2562 2817 2568
rect 2886 2562 2889 2588
rect 2926 2582 2929 2658
rect 2942 2612 2945 2668
rect 2966 2622 2969 2658
rect 2894 2552 2897 2568
rect 2874 2548 2878 2551
rect 2818 2538 2822 2541
rect 2842 2538 2846 2541
rect 2838 2522 2841 2528
rect 2814 2462 2817 2468
rect 2782 2452 2785 2458
rect 2818 2448 2822 2451
rect 2790 2442 2793 2448
rect 2806 2442 2809 2448
rect 2830 2402 2833 2458
rect 2838 2442 2841 2518
rect 2862 2502 2865 2538
rect 2846 2492 2849 2498
rect 2886 2492 2889 2518
rect 2902 2472 2905 2518
rect 2918 2492 2921 2558
rect 2934 2552 2937 2598
rect 2958 2572 2961 2578
rect 2966 2551 2969 2608
rect 2962 2548 2969 2551
rect 2942 2501 2945 2538
rect 2950 2512 2953 2538
rect 2938 2498 2945 2501
rect 2854 2452 2857 2468
rect 2898 2458 2902 2461
rect 2918 2452 2921 2488
rect 2934 2472 2937 2498
rect 2966 2462 2969 2468
rect 2946 2458 2950 2461
rect 2954 2448 2958 2451
rect 2718 2352 2721 2388
rect 2786 2368 2790 2371
rect 2746 2358 2750 2361
rect 2818 2358 2822 2361
rect 2682 2348 2686 2351
rect 2738 2348 2742 2351
rect 2670 2338 2678 2341
rect 2694 2332 2697 2348
rect 2594 2328 2598 2331
rect 2666 2328 2670 2331
rect 2646 2311 2649 2318
rect 2646 2308 2657 2311
rect 2494 2242 2497 2258
rect 2462 2152 2465 2158
rect 2502 2152 2505 2278
rect 2582 2272 2585 2298
rect 2590 2292 2593 2298
rect 2646 2292 2649 2298
rect 2602 2278 2606 2281
rect 2574 2262 2577 2268
rect 2518 2212 2521 2258
rect 2536 2203 2538 2207
rect 2542 2203 2545 2207
rect 2549 2203 2552 2207
rect 2518 2162 2521 2168
rect 2390 2142 2393 2148
rect 2414 2132 2417 2138
rect 2278 2092 2281 2108
rect 2290 2078 2294 2081
rect 2306 2078 2310 2081
rect 2326 2072 2329 2108
rect 2334 2072 2337 2118
rect 2350 2102 2353 2118
rect 2394 2078 2401 2081
rect 2410 2078 2414 2081
rect 2382 2072 2385 2078
rect 2398 2072 2401 2078
rect 2290 2068 2294 2071
rect 2318 2062 2321 2068
rect 2422 2062 2425 2118
rect 2430 2072 2433 2128
rect 2442 2078 2446 2081
rect 2454 2081 2457 2128
rect 2450 2078 2457 2081
rect 2462 2071 2465 2118
rect 2486 2082 2489 2128
rect 2458 2068 2465 2071
rect 2394 2058 2398 2061
rect 2254 1982 2257 2018
rect 2270 1992 2273 2058
rect 2302 2052 2305 2058
rect 2110 1962 2113 1968
rect 2146 1958 2150 1961
rect 2178 1958 2182 1961
rect 2062 1892 2065 1908
rect 2094 1892 2097 1918
rect 2078 1852 2081 1858
rect 2086 1802 2089 1868
rect 1998 1752 2001 1778
rect 1990 1672 1993 1728
rect 1998 1662 2001 1708
rect 2006 1681 2009 1768
rect 2042 1748 2046 1751
rect 2042 1738 2046 1741
rect 2030 1722 2033 1728
rect 2024 1703 2026 1707
rect 2030 1703 2033 1707
rect 2037 1703 2040 1707
rect 2054 1702 2057 1758
rect 2062 1752 2065 1758
rect 2078 1752 2081 1798
rect 2086 1742 2089 1798
rect 2094 1772 2097 1838
rect 2062 1682 2065 1688
rect 2006 1678 2014 1681
rect 1982 1652 1985 1658
rect 2018 1568 2022 1571
rect 1890 1528 1894 1531
rect 1878 1518 1889 1521
rect 1886 1492 1889 1518
rect 1902 1482 1905 1538
rect 1910 1502 1913 1548
rect 1918 1532 1921 1538
rect 1934 1492 1937 1548
rect 1942 1532 1945 1558
rect 1950 1548 1958 1551
rect 1950 1521 1953 1548
rect 1966 1542 1969 1548
rect 1942 1518 1953 1521
rect 1902 1472 1905 1478
rect 1862 1462 1865 1468
rect 1854 1342 1857 1428
rect 1870 1412 1873 1468
rect 1878 1432 1881 1468
rect 1902 1458 1910 1461
rect 1914 1458 1918 1461
rect 1886 1448 1894 1451
rect 1886 1372 1889 1448
rect 1902 1382 1905 1458
rect 1926 1442 1929 1448
rect 1910 1362 1913 1418
rect 1918 1412 1921 1438
rect 1934 1412 1937 1448
rect 1918 1392 1921 1398
rect 1942 1372 1945 1518
rect 1974 1512 1977 1548
rect 1982 1528 1990 1531
rect 1986 1518 1990 1521
rect 1950 1462 1953 1508
rect 1990 1492 1993 1508
rect 1998 1482 2001 1558
rect 2006 1551 2009 1568
rect 2030 1552 2033 1568
rect 2006 1548 2014 1551
rect 2022 1542 2025 1548
rect 2038 1532 2041 1658
rect 2014 1528 2022 1531
rect 2014 1502 2017 1528
rect 2024 1503 2026 1507
rect 2030 1503 2033 1507
rect 2037 1503 2040 1507
rect 2046 1492 2049 1648
rect 2054 1562 2057 1678
rect 2070 1592 2073 1738
rect 2078 1712 2081 1728
rect 2094 1711 2097 1768
rect 2102 1762 2105 1918
rect 2118 1912 2121 1948
rect 2166 1942 2169 1948
rect 2130 1938 2134 1941
rect 2146 1928 2150 1931
rect 2118 1882 2121 1908
rect 2134 1902 2137 1928
rect 2158 1912 2161 1938
rect 2182 1882 2185 1928
rect 2190 1892 2193 1908
rect 2198 1902 2201 1948
rect 2206 1912 2209 1978
rect 2262 1962 2265 1968
rect 2230 1952 2233 1958
rect 2218 1928 2222 1931
rect 2206 1882 2209 1908
rect 2214 1892 2217 1898
rect 2138 1868 2142 1871
rect 2170 1868 2174 1871
rect 2118 1862 2121 1868
rect 2110 1851 2113 1858
rect 2110 1848 2121 1851
rect 2110 1792 2113 1798
rect 2118 1772 2121 1848
rect 2122 1758 2126 1761
rect 2142 1752 2145 1858
rect 2150 1802 2153 1868
rect 2150 1792 2153 1798
rect 2158 1792 2161 1858
rect 2178 1848 2185 1851
rect 2122 1748 2126 1751
rect 2154 1748 2169 1751
rect 2102 1742 2105 1748
rect 2166 1742 2169 1748
rect 2154 1738 2158 1741
rect 2106 1728 2110 1731
rect 2086 1708 2097 1711
rect 2086 1682 2089 1708
rect 2118 1702 2121 1728
rect 2126 1712 2129 1738
rect 2142 1731 2145 1738
rect 2142 1728 2150 1731
rect 2166 1712 2169 1728
rect 2174 1722 2177 1748
rect 2182 1742 2185 1848
rect 2190 1762 2193 1788
rect 2198 1752 2201 1868
rect 2206 1862 2209 1878
rect 2230 1872 2233 1938
rect 2238 1932 2241 1938
rect 2246 1912 2249 1948
rect 2270 1932 2273 1948
rect 2254 1892 2257 1928
rect 2278 1892 2281 1958
rect 2286 1932 2289 2038
rect 2294 1942 2297 2018
rect 2318 1952 2321 1958
rect 2350 1952 2353 2048
rect 2366 2042 2369 2048
rect 2382 1992 2385 2058
rect 2430 2052 2433 2068
rect 2462 2052 2465 2058
rect 2486 2052 2489 2068
rect 2414 2042 2417 2048
rect 2478 2042 2481 2048
rect 2450 2038 2454 2041
rect 2370 1958 2374 1961
rect 2394 1958 2398 1961
rect 2406 1952 2409 2038
rect 2386 1948 2390 1951
rect 2338 1938 2342 1941
rect 2294 1932 2297 1938
rect 2238 1882 2241 1888
rect 2246 1882 2249 1888
rect 2294 1872 2297 1888
rect 2310 1881 2313 1918
rect 2318 1892 2321 1938
rect 2330 1928 2334 1931
rect 2326 1892 2329 1918
rect 2350 1882 2353 1948
rect 2310 1878 2321 1881
rect 2234 1868 2238 1871
rect 2254 1868 2262 1871
rect 2254 1792 2257 1868
rect 2270 1852 2273 1858
rect 2278 1852 2281 1858
rect 2198 1722 2201 1738
rect 2174 1712 2177 1718
rect 2094 1692 2097 1698
rect 2134 1692 2137 1698
rect 2198 1692 2201 1698
rect 2162 1688 2166 1691
rect 2078 1672 2081 1678
rect 2126 1672 2129 1688
rect 2078 1652 2081 1658
rect 2082 1648 2089 1651
rect 2086 1552 2089 1648
rect 2094 1552 2097 1558
rect 2078 1512 2081 1548
rect 2090 1528 2094 1531
rect 2102 1521 2105 1668
rect 2110 1652 2113 1658
rect 2118 1652 2121 1658
rect 2142 1622 2145 1678
rect 2150 1622 2153 1688
rect 2206 1682 2209 1758
rect 2222 1752 2225 1778
rect 2214 1742 2217 1748
rect 2230 1732 2233 1758
rect 2254 1742 2257 1748
rect 2230 1682 2233 1688
rect 2186 1668 2190 1671
rect 2166 1662 2169 1668
rect 2214 1662 2217 1678
rect 2238 1671 2241 1678
rect 2262 1672 2265 1828
rect 2270 1792 2273 1848
rect 2270 1742 2273 1758
rect 2282 1748 2286 1751
rect 2294 1741 2297 1858
rect 2302 1852 2305 1858
rect 2310 1812 2313 1868
rect 2310 1792 2313 1808
rect 2286 1738 2297 1741
rect 2302 1742 2305 1758
rect 2318 1752 2321 1878
rect 2326 1852 2329 1878
rect 2334 1872 2337 1878
rect 2358 1872 2361 1948
rect 2366 1938 2374 1941
rect 2346 1868 2350 1871
rect 2334 1812 2337 1868
rect 2366 1862 2369 1938
rect 2334 1782 2337 1788
rect 2278 1702 2281 1738
rect 2286 1692 2289 1738
rect 2306 1728 2310 1731
rect 2318 1692 2321 1728
rect 2342 1721 2345 1828
rect 2366 1752 2369 1778
rect 2334 1718 2345 1721
rect 2334 1682 2337 1718
rect 2342 1692 2345 1708
rect 2350 1692 2353 1748
rect 2358 1732 2361 1738
rect 2274 1678 2278 1681
rect 2366 1672 2369 1698
rect 2374 1692 2377 1918
rect 2406 1892 2409 1948
rect 2390 1782 2393 1868
rect 2414 1831 2417 2008
rect 2422 1992 2425 1998
rect 2446 1992 2449 2008
rect 2466 1988 2470 1991
rect 2462 1952 2465 1978
rect 2478 1942 2481 2028
rect 2494 2012 2497 2138
rect 2502 2092 2505 2138
rect 2526 2132 2529 2138
rect 2510 2082 2513 2098
rect 2518 2082 2521 2118
rect 2534 2102 2537 2118
rect 2542 2082 2545 2168
rect 2558 2152 2561 2218
rect 2554 2078 2558 2081
rect 2502 2071 2505 2078
rect 2502 2068 2513 2071
rect 2486 1952 2489 1958
rect 2502 1932 2505 2018
rect 2494 1912 2497 1918
rect 2454 1892 2457 1908
rect 2494 1892 2497 1898
rect 2510 1892 2513 2068
rect 2534 2022 2537 2068
rect 2518 2012 2521 2018
rect 2536 2003 2538 2007
rect 2542 2003 2545 2007
rect 2549 2003 2552 2007
rect 2518 1992 2521 1998
rect 2558 1991 2561 2008
rect 2550 1988 2561 1991
rect 2566 1992 2569 2198
rect 2574 2192 2577 2258
rect 2606 2252 2609 2258
rect 2598 2152 2601 2158
rect 2622 2152 2625 2288
rect 2634 2268 2638 2271
rect 2638 2242 2641 2248
rect 2654 2172 2657 2308
rect 2678 2282 2681 2298
rect 2710 2292 2713 2318
rect 2726 2312 2729 2338
rect 2662 2262 2665 2278
rect 2686 2272 2689 2288
rect 2702 2272 2705 2278
rect 2734 2272 2737 2278
rect 2698 2258 2702 2261
rect 2706 2258 2710 2261
rect 2658 2148 2662 2151
rect 2550 1952 2553 1988
rect 2582 1962 2585 2118
rect 2590 2042 2593 2048
rect 2598 2022 2601 2148
rect 2606 2142 2609 2148
rect 2606 2092 2609 2098
rect 2610 2068 2614 2071
rect 2622 2061 2625 2148
rect 2630 2142 2633 2148
rect 2678 2141 2681 2258
rect 2718 2252 2721 2258
rect 2734 2252 2737 2258
rect 2742 2252 2745 2268
rect 2750 2262 2753 2328
rect 2758 2282 2761 2338
rect 2806 2332 2809 2338
rect 2782 2292 2785 2298
rect 2814 2291 2817 2358
rect 2830 2352 2833 2368
rect 2846 2341 2849 2418
rect 2842 2338 2849 2341
rect 2822 2312 2825 2338
rect 2814 2288 2825 2291
rect 2802 2278 2806 2281
rect 2766 2272 2769 2278
rect 2814 2272 2817 2278
rect 2758 2262 2761 2268
rect 2766 2262 2769 2268
rect 2754 2258 2758 2261
rect 2706 2248 2710 2251
rect 2718 2182 2721 2248
rect 2742 2242 2745 2248
rect 2758 2192 2761 2218
rect 2690 2148 2694 2151
rect 2702 2142 2705 2148
rect 2726 2142 2729 2158
rect 2746 2148 2750 2151
rect 2766 2142 2769 2248
rect 2774 2212 2777 2248
rect 2798 2192 2801 2208
rect 2814 2202 2817 2258
rect 2822 2252 2825 2288
rect 2838 2262 2841 2328
rect 2846 2272 2849 2338
rect 2854 2312 2857 2448
rect 2870 2392 2873 2438
rect 2890 2418 2894 2421
rect 2862 2332 2865 2358
rect 2870 2352 2873 2368
rect 2918 2362 2921 2448
rect 2966 2442 2969 2448
rect 2974 2412 2977 2668
rect 3022 2661 3025 2708
rect 3030 2672 3033 2728
rect 3038 2722 3041 2758
rect 3054 2732 3057 2838
rect 3070 2752 3073 2758
rect 3078 2742 3081 2878
rect 3086 2852 3089 2858
rect 3094 2842 3097 2928
rect 3102 2872 3105 2878
rect 3110 2871 3113 2948
rect 3118 2892 3121 2948
rect 3130 2938 3134 2941
rect 3154 2938 3158 2941
rect 3142 2932 3145 2938
rect 3174 2932 3177 2948
rect 3126 2922 3129 2928
rect 3158 2922 3161 2928
rect 3118 2872 3121 2878
rect 3110 2868 3118 2871
rect 3110 2842 3113 2848
rect 3086 2752 3089 2788
rect 3086 2742 3089 2748
rect 3040 2703 3042 2707
rect 3046 2703 3049 2707
rect 3053 2703 3056 2707
rect 3042 2688 3046 2691
rect 3078 2672 3081 2738
rect 3094 2732 3097 2818
rect 3110 2742 3113 2768
rect 3102 2711 3105 2718
rect 3102 2708 3113 2711
rect 3102 2662 3105 2698
rect 3022 2658 3030 2661
rect 2982 2652 2985 2658
rect 2998 2652 3001 2658
rect 2982 2562 2985 2648
rect 3006 2592 3009 2618
rect 3014 2552 3017 2568
rect 2998 2522 3001 2548
rect 3006 2542 3009 2548
rect 3022 2532 3025 2538
rect 3038 2532 3041 2588
rect 3050 2568 3054 2571
rect 3070 2562 3073 2658
rect 3078 2552 3081 2578
rect 2998 2482 3001 2518
rect 2990 2472 2993 2478
rect 3014 2472 3017 2508
rect 3030 2492 3033 2518
rect 3040 2503 3042 2507
rect 3046 2503 3049 2507
rect 3053 2503 3056 2507
rect 3062 2482 3065 2528
rect 3026 2458 3030 2461
rect 2982 2452 2985 2458
rect 3014 2451 3017 2458
rect 3038 2452 3041 2468
rect 3014 2448 3022 2451
rect 3062 2442 3065 2478
rect 3074 2468 3078 2471
rect 3086 2461 3089 2648
rect 3110 2591 3113 2708
rect 3118 2672 3121 2738
rect 3118 2642 3121 2668
rect 3110 2588 3121 2591
rect 3098 2558 3102 2561
rect 3094 2542 3097 2558
rect 3110 2542 3113 2578
rect 3118 2562 3121 2588
rect 3126 2542 3129 2868
rect 3150 2812 3153 2848
rect 3158 2812 3161 2918
rect 3182 2912 3185 2958
rect 3262 2952 3265 2958
rect 3278 2952 3281 2958
rect 3334 2952 3337 3038
rect 3226 2948 3230 2951
rect 3306 2948 3310 2951
rect 3190 2942 3193 2948
rect 3198 2922 3201 2948
rect 3206 2932 3209 2938
rect 3214 2912 3217 2938
rect 3246 2912 3249 2948
rect 3254 2942 3257 2948
rect 3294 2932 3297 2938
rect 3274 2928 3278 2931
rect 3186 2878 3190 2881
rect 3182 2862 3185 2868
rect 3190 2862 3193 2878
rect 3206 2872 3209 2878
rect 3214 2871 3217 2908
rect 3254 2892 3257 2928
rect 3234 2878 3238 2881
rect 3214 2868 3222 2871
rect 3202 2858 3206 2861
rect 3174 2822 3177 2828
rect 3138 2758 3142 2761
rect 3138 2748 3142 2751
rect 3134 2692 3137 2728
rect 3134 2662 3137 2668
rect 3134 2552 3137 2648
rect 3142 2592 3145 2718
rect 3158 2712 3161 2748
rect 3166 2742 3169 2758
rect 3174 2742 3177 2808
rect 3194 2758 3198 2761
rect 3182 2752 3185 2758
rect 3174 2731 3177 2738
rect 3166 2728 3177 2731
rect 3190 2732 3193 2738
rect 3198 2732 3201 2758
rect 3206 2732 3209 2818
rect 3214 2812 3217 2858
rect 3222 2772 3225 2868
rect 3246 2862 3249 2868
rect 3262 2862 3265 2878
rect 3270 2872 3273 2918
rect 3254 2858 3262 2861
rect 3238 2762 3241 2818
rect 3234 2748 3238 2751
rect 3150 2672 3153 2698
rect 3166 2692 3169 2728
rect 3174 2682 3177 2698
rect 3198 2682 3201 2718
rect 3206 2682 3209 2688
rect 3182 2662 3185 2668
rect 3198 2662 3201 2668
rect 3154 2658 3158 2661
rect 3150 2552 3153 2638
rect 3182 2562 3185 2618
rect 3198 2582 3201 2658
rect 3206 2602 3209 2678
rect 3198 2552 3201 2568
rect 3206 2542 3209 2598
rect 3154 2538 3158 2541
rect 3142 2532 3145 2538
rect 3170 2528 3174 2531
rect 3182 2522 3185 2528
rect 3078 2458 3089 2461
rect 3078 2452 3081 2458
rect 2934 2372 2937 2378
rect 2950 2362 2953 2368
rect 2962 2358 2966 2361
rect 2906 2348 2910 2351
rect 2938 2348 2942 2351
rect 2954 2348 2958 2351
rect 2870 2332 2873 2348
rect 2930 2338 2934 2341
rect 2886 2332 2889 2338
rect 2866 2318 2870 2321
rect 2918 2312 2921 2328
rect 2854 2272 2857 2288
rect 2838 2222 2841 2258
rect 2806 2162 2809 2168
rect 2822 2162 2825 2168
rect 2834 2158 2838 2161
rect 2774 2152 2777 2158
rect 2826 2148 2830 2151
rect 2782 2142 2785 2148
rect 2678 2138 2686 2141
rect 2670 2132 2673 2138
rect 2630 2092 2633 2128
rect 2646 2112 2649 2118
rect 2678 2091 2681 2118
rect 2670 2088 2681 2091
rect 2670 2072 2673 2088
rect 2678 2072 2681 2078
rect 2614 2058 2625 2061
rect 2674 2058 2678 2061
rect 2554 1938 2558 1941
rect 2566 1932 2569 1948
rect 2590 1932 2593 2018
rect 2606 1952 2609 1958
rect 2614 1952 2617 2058
rect 2646 1952 2649 2058
rect 2686 2052 2689 2138
rect 2694 2132 2697 2138
rect 2702 2052 2705 2138
rect 2718 2102 2721 2128
rect 2726 2092 2729 2138
rect 2742 2102 2745 2138
rect 2794 2128 2798 2131
rect 2714 2088 2718 2091
rect 2734 2072 2737 2078
rect 2742 2052 2745 2098
rect 2750 2052 2753 2108
rect 2758 2072 2761 2078
rect 2758 2052 2761 2068
rect 2766 2062 2769 2078
rect 2782 2072 2785 2078
rect 2790 2062 2793 2088
rect 2798 2062 2801 2098
rect 2814 2052 2817 2078
rect 2654 2042 2657 2048
rect 2718 2042 2721 2048
rect 2750 2042 2753 2048
rect 2762 2038 2766 2041
rect 2678 1952 2681 1958
rect 2650 1948 2654 1951
rect 2450 1868 2454 1871
rect 2430 1842 2433 1868
rect 2486 1852 2489 1868
rect 2526 1862 2529 1868
rect 2574 1862 2577 1908
rect 2590 1852 2593 1878
rect 2414 1828 2425 1831
rect 2414 1812 2417 1818
rect 2414 1752 2417 1798
rect 2390 1732 2393 1748
rect 2382 1702 2385 1718
rect 2230 1668 2241 1671
rect 2174 1641 2177 1658
rect 2182 1652 2185 1658
rect 2222 1651 2225 1668
rect 2214 1648 2225 1651
rect 2174 1638 2185 1641
rect 2146 1578 2150 1581
rect 2134 1562 2137 1578
rect 2182 1572 2185 1638
rect 2214 1592 2217 1648
rect 2230 1572 2233 1668
rect 2246 1651 2249 1668
rect 2254 1662 2257 1668
rect 2246 1648 2257 1651
rect 2238 1592 2241 1608
rect 2254 1592 2257 1648
rect 2270 1642 2273 1648
rect 2218 1568 2225 1571
rect 2086 1518 2105 1521
rect 2154 1548 2158 1551
rect 2110 1542 2113 1548
rect 2110 1522 2113 1538
rect 2086 1501 2089 1518
rect 2118 1502 2121 1548
rect 2126 1542 2129 1548
rect 2134 1512 2137 1548
rect 2174 1542 2177 1568
rect 2190 1552 2193 1558
rect 2190 1542 2193 1548
rect 2214 1532 2217 1548
rect 2222 1542 2225 1568
rect 2254 1561 2257 1578
rect 2254 1558 2262 1561
rect 2266 1538 2270 1541
rect 2078 1498 2089 1501
rect 2078 1492 2081 1498
rect 2102 1492 2105 1498
rect 2166 1492 2169 1498
rect 1958 1442 1961 1468
rect 1966 1462 1969 1478
rect 1982 1441 1985 1478
rect 2046 1472 2049 1488
rect 2002 1458 2006 1461
rect 1990 1442 1993 1448
rect 1982 1438 1990 1441
rect 1958 1432 1961 1438
rect 1950 1412 1953 1418
rect 1874 1358 1878 1361
rect 1898 1358 1902 1361
rect 1942 1352 1945 1358
rect 1914 1348 1918 1351
rect 1902 1342 1905 1348
rect 1918 1332 1921 1338
rect 1934 1332 1937 1338
rect 1842 1328 1846 1331
rect 1882 1328 1886 1331
rect 1886 1312 1889 1328
rect 1942 1322 1945 1338
rect 1854 1292 1857 1298
rect 1794 1268 1798 1271
rect 1774 1238 1785 1241
rect 1746 1228 1750 1231
rect 1686 1152 1689 1158
rect 1694 1152 1697 1158
rect 1750 1152 1753 1158
rect 1758 1152 1761 1178
rect 1774 1162 1777 1238
rect 1794 1188 1798 1191
rect 1730 1148 1734 1151
rect 1706 1138 1710 1141
rect 1730 1138 1734 1141
rect 1742 1131 1745 1148
rect 1750 1142 1753 1148
rect 1734 1128 1745 1131
rect 1686 1082 1689 1088
rect 1694 1072 1697 1118
rect 1670 1052 1673 1058
rect 1650 1048 1654 1051
rect 1630 1038 1641 1041
rect 1630 942 1633 1038
rect 1670 992 1673 1008
rect 1678 1002 1681 1068
rect 1702 1052 1705 1128
rect 1718 1102 1721 1128
rect 1734 1092 1737 1128
rect 1750 1082 1753 1128
rect 1726 1072 1729 1078
rect 1714 1068 1718 1071
rect 1686 1012 1689 1048
rect 1694 1042 1697 1048
rect 1710 1042 1713 1048
rect 1718 1012 1721 1058
rect 1734 1012 1737 1078
rect 1742 1052 1745 1078
rect 1758 1062 1761 1138
rect 1766 1082 1769 1158
rect 1774 1152 1777 1158
rect 1806 1152 1809 1288
rect 1822 1278 1830 1281
rect 1878 1281 1881 1308
rect 1894 1292 1897 1308
rect 1910 1281 1913 1298
rect 1878 1278 1889 1281
rect 1910 1278 1921 1281
rect 1822 1272 1825 1278
rect 1846 1272 1849 1278
rect 1834 1268 1838 1271
rect 1870 1262 1873 1278
rect 1878 1262 1881 1268
rect 1818 1258 1822 1261
rect 1886 1252 1889 1278
rect 1906 1268 1910 1271
rect 1918 1262 1921 1278
rect 1906 1258 1913 1261
rect 1838 1248 1846 1251
rect 1894 1251 1897 1258
rect 1926 1251 1929 1288
rect 1934 1262 1937 1308
rect 1950 1302 1953 1368
rect 1958 1352 1961 1428
rect 1950 1272 1953 1288
rect 1966 1282 1969 1418
rect 1974 1372 1977 1418
rect 1998 1412 2001 1428
rect 1974 1352 1977 1358
rect 1982 1342 1985 1348
rect 1990 1332 1993 1338
rect 1974 1282 1977 1298
rect 1894 1248 1929 1251
rect 1942 1251 1945 1268
rect 1950 1262 1953 1268
rect 1938 1248 1945 1251
rect 1814 1232 1817 1238
rect 1822 1162 1825 1248
rect 1830 1212 1833 1228
rect 1838 1212 1841 1248
rect 1990 1232 1993 1318
rect 1998 1272 2001 1318
rect 2006 1272 2009 1448
rect 2014 1382 2017 1468
rect 2074 1458 2078 1461
rect 2070 1432 2073 1448
rect 2086 1442 2089 1468
rect 2094 1452 2097 1478
rect 2122 1468 2126 1471
rect 2014 1332 2017 1358
rect 2046 1342 2049 1368
rect 2058 1348 2062 1351
rect 2070 1351 2073 1388
rect 2070 1348 2081 1351
rect 2062 1332 2065 1338
rect 2038 1322 2041 1328
rect 2070 1322 2073 1338
rect 2078 1332 2081 1348
rect 2086 1342 2089 1398
rect 2102 1382 2105 1468
rect 2110 1462 2113 1468
rect 2150 1462 2153 1468
rect 2130 1458 2134 1461
rect 2118 1452 2121 1458
rect 2146 1448 2150 1451
rect 2102 1362 2105 1368
rect 2110 1362 2113 1408
rect 2098 1348 2102 1351
rect 2110 1341 2113 1348
rect 2102 1338 2113 1341
rect 2118 1342 2121 1368
rect 2150 1342 2153 1388
rect 2158 1352 2161 1478
rect 2178 1468 2182 1471
rect 2174 1452 2177 1458
rect 2174 1352 2177 1398
rect 2182 1392 2185 1448
rect 2190 1362 2193 1488
rect 2206 1472 2209 1488
rect 2214 1472 2217 1478
rect 2222 1462 2225 1538
rect 2230 1502 2233 1538
rect 2278 1532 2281 1628
rect 2286 1552 2289 1658
rect 2294 1652 2297 1668
rect 2302 1632 2305 1658
rect 2310 1632 2313 1668
rect 2326 1602 2329 1648
rect 2334 1628 2342 1631
rect 2306 1588 2310 1591
rect 2306 1558 2310 1561
rect 2314 1538 2318 1541
rect 2286 1532 2289 1538
rect 2242 1528 2246 1531
rect 2270 1478 2278 1481
rect 2218 1458 2222 1461
rect 2242 1458 2246 1461
rect 2198 1452 2201 1458
rect 2024 1303 2026 1307
rect 2030 1303 2033 1307
rect 2037 1303 2040 1307
rect 2078 1282 2081 1318
rect 2086 1282 2089 1298
rect 2094 1282 2097 1328
rect 2102 1292 2105 1338
rect 2130 1328 2134 1331
rect 2110 1322 2113 1328
rect 2034 1278 2038 1281
rect 2086 1272 2089 1278
rect 2046 1268 2081 1271
rect 1970 1218 1974 1221
rect 1838 1202 1841 1208
rect 1858 1188 1862 1191
rect 1802 1138 1806 1141
rect 1774 1102 1777 1138
rect 1814 1131 1817 1158
rect 1830 1152 1833 1158
rect 1846 1142 1849 1188
rect 1858 1148 1862 1151
rect 1870 1141 1873 1148
rect 1850 1138 1857 1141
rect 1806 1128 1817 1131
rect 1834 1128 1838 1131
rect 1782 1081 1785 1128
rect 1790 1092 1793 1128
rect 1806 1082 1809 1128
rect 1814 1102 1817 1118
rect 1830 1082 1833 1118
rect 1838 1082 1841 1088
rect 1782 1078 1793 1081
rect 1802 1078 1806 1081
rect 1774 1062 1777 1078
rect 1790 1072 1793 1078
rect 1846 1071 1849 1078
rect 1842 1068 1849 1071
rect 1766 1051 1769 1058
rect 1762 1048 1769 1051
rect 1734 992 1737 1008
rect 1742 992 1745 1008
rect 1646 962 1649 968
rect 1718 952 1721 958
rect 1750 952 1753 958
rect 1682 948 1686 951
rect 1694 942 1697 948
rect 1718 942 1721 948
rect 1582 872 1585 938
rect 1590 872 1593 898
rect 1446 852 1449 858
rect 1478 852 1481 858
rect 1430 841 1433 848
rect 1414 838 1433 841
rect 1310 798 1318 801
rect 1310 792 1313 798
rect 1366 792 1369 808
rect 1406 792 1409 808
rect 1454 792 1457 838
rect 1462 812 1465 848
rect 1266 738 1273 741
rect 1254 721 1257 728
rect 1246 718 1257 721
rect 1230 681 1233 698
rect 1246 692 1249 718
rect 1270 692 1273 738
rect 1294 712 1297 748
rect 1302 742 1305 748
rect 1310 732 1313 778
rect 1334 771 1337 778
rect 1334 768 1350 771
rect 1394 768 1398 771
rect 1414 762 1417 768
rect 1334 742 1337 748
rect 1326 732 1329 738
rect 1342 692 1345 748
rect 1350 742 1353 748
rect 1374 732 1377 748
rect 1406 742 1409 748
rect 1422 742 1425 748
rect 1230 678 1238 681
rect 1362 678 1366 681
rect 1206 672 1209 678
rect 1174 622 1177 648
rect 1198 582 1201 668
rect 1214 662 1217 678
rect 1262 672 1265 678
rect 1310 672 1313 678
rect 1334 672 1337 678
rect 1390 672 1393 678
rect 1290 668 1294 671
rect 1254 662 1257 668
rect 1274 658 1278 661
rect 1298 658 1302 661
rect 1214 632 1217 638
rect 1222 632 1225 658
rect 1230 652 1233 658
rect 1206 592 1209 628
rect 1238 612 1241 648
rect 1286 642 1289 648
rect 1198 572 1201 578
rect 1310 571 1313 668
rect 1322 658 1326 661
rect 1334 582 1337 658
rect 1366 652 1369 658
rect 1346 638 1350 641
rect 1342 592 1345 608
rect 1310 568 1318 571
rect 1326 568 1334 571
rect 1294 562 1297 568
rect 1226 558 1230 561
rect 1286 552 1289 558
rect 1194 548 1198 551
rect 1182 542 1185 548
rect 1198 532 1201 538
rect 1206 502 1209 548
rect 1222 492 1225 528
rect 1246 512 1249 548
rect 1270 522 1273 528
rect 1270 492 1273 498
rect 1142 462 1145 468
rect 1190 462 1193 468
rect 1206 462 1209 468
rect 1230 462 1233 468
rect 1310 462 1313 548
rect 1318 542 1321 548
rect 1326 522 1329 568
rect 1334 558 1342 561
rect 1318 492 1321 508
rect 1326 462 1329 468
rect 1114 458 1118 461
rect 1282 458 1286 461
rect 1094 452 1097 458
rect 1062 378 1073 381
rect 1026 348 1030 351
rect 1030 292 1033 318
rect 1022 282 1025 288
rect 1038 272 1041 278
rect 1054 271 1057 348
rect 1062 292 1065 378
rect 1070 352 1073 358
rect 1046 268 1057 271
rect 926 222 929 258
rect 934 242 937 268
rect 950 262 953 268
rect 1046 262 1049 268
rect 990 252 993 258
rect 1038 252 1041 258
rect 870 112 873 138
rect 910 112 913 178
rect 834 68 838 71
rect 806 62 809 68
rect 702 32 705 38
rect 782 32 785 48
rect 790 42 793 48
rect 814 42 817 68
rect 822 62 825 68
rect 862 52 865 98
rect 886 92 889 98
rect 870 62 873 68
rect 910 61 913 108
rect 918 92 921 168
rect 934 161 937 238
rect 966 192 969 248
rect 1046 242 1049 258
rect 930 158 937 161
rect 926 142 929 158
rect 950 152 953 158
rect 954 138 958 141
rect 982 132 985 158
rect 998 142 1001 198
rect 1030 192 1033 198
rect 1046 142 1049 178
rect 1054 152 1057 258
rect 1070 192 1073 288
rect 1086 251 1089 378
rect 1094 322 1097 348
rect 1094 292 1097 318
rect 1102 282 1105 458
rect 1126 392 1129 398
rect 1134 392 1137 458
rect 1150 422 1153 458
rect 1158 452 1161 458
rect 1170 418 1177 421
rect 1174 392 1177 418
rect 1110 352 1113 358
rect 1138 348 1142 351
rect 1154 348 1158 351
rect 1170 348 1174 351
rect 1118 322 1121 348
rect 1110 272 1113 278
rect 1082 248 1089 251
rect 1094 242 1097 258
rect 1102 252 1105 268
rect 1118 262 1121 298
rect 1142 282 1145 288
rect 1126 278 1134 281
rect 1126 272 1129 278
rect 1166 272 1169 278
rect 1174 272 1177 338
rect 1182 302 1185 458
rect 1198 382 1201 458
rect 1230 392 1233 458
rect 1246 432 1249 458
rect 1254 452 1257 458
rect 1294 432 1297 458
rect 1302 392 1305 458
rect 1254 352 1257 358
rect 1286 352 1289 358
rect 1326 352 1329 408
rect 1334 382 1337 558
rect 1358 552 1361 628
rect 1374 592 1377 648
rect 1382 582 1385 618
rect 1366 552 1369 558
rect 1390 552 1393 658
rect 1398 652 1401 698
rect 1430 681 1433 778
rect 1478 772 1481 788
rect 1486 772 1489 868
rect 1494 842 1497 858
rect 1502 792 1505 818
rect 1512 803 1514 807
rect 1518 803 1521 807
rect 1525 803 1528 807
rect 1522 788 1526 791
rect 1534 772 1537 868
rect 1542 812 1545 868
rect 1578 858 1582 861
rect 1586 848 1590 851
rect 1554 838 1558 841
rect 1566 832 1569 848
rect 1570 768 1574 771
rect 1486 762 1489 768
rect 1438 712 1441 728
rect 1422 678 1433 681
rect 1422 672 1425 678
rect 1410 658 1414 661
rect 1430 652 1433 668
rect 1446 661 1449 758
rect 1590 752 1593 758
rect 1442 658 1449 661
rect 1462 662 1465 738
rect 1470 722 1473 728
rect 1470 682 1473 688
rect 1478 672 1481 728
rect 1474 668 1478 671
rect 1486 671 1489 748
rect 1550 742 1553 748
rect 1590 742 1593 748
rect 1566 738 1574 741
rect 1514 728 1518 731
rect 1502 722 1505 728
rect 1514 678 1518 681
rect 1486 668 1494 671
rect 1494 662 1497 668
rect 1414 602 1417 618
rect 1386 548 1390 551
rect 1342 542 1345 548
rect 1358 512 1361 548
rect 1342 472 1345 508
rect 1406 492 1409 548
rect 1414 542 1417 548
rect 1438 532 1441 548
rect 1426 518 1430 521
rect 1430 492 1433 498
rect 1438 492 1441 498
rect 1430 482 1433 488
rect 1446 472 1449 658
rect 1458 648 1462 651
rect 1478 592 1481 648
rect 1486 632 1489 658
rect 1482 548 1486 551
rect 1454 542 1457 548
rect 1462 512 1465 548
rect 1342 392 1345 458
rect 1374 402 1377 418
rect 1390 412 1393 468
rect 1398 462 1401 468
rect 1410 458 1414 461
rect 1422 452 1425 468
rect 1478 462 1481 508
rect 1494 492 1497 658
rect 1502 648 1510 651
rect 1502 572 1505 648
rect 1512 603 1514 607
rect 1518 603 1521 607
rect 1525 603 1528 607
rect 1534 592 1537 658
rect 1518 552 1521 558
rect 1526 532 1529 548
rect 1522 468 1526 471
rect 1430 452 1433 458
rect 1446 422 1449 458
rect 1430 392 1433 418
rect 1398 352 1401 388
rect 1430 372 1433 388
rect 1210 348 1214 351
rect 1234 348 1238 351
rect 1354 348 1358 351
rect 1190 292 1193 348
rect 1198 322 1201 348
rect 1154 258 1158 261
rect 1174 258 1182 261
rect 1118 252 1121 258
rect 1166 251 1169 258
rect 1146 248 1169 251
rect 1126 192 1129 228
rect 1174 192 1177 258
rect 1190 232 1193 248
rect 1198 242 1201 318
rect 1222 292 1225 348
rect 1266 338 1270 341
rect 1238 262 1241 338
rect 1278 322 1281 348
rect 1246 292 1249 308
rect 1254 302 1257 308
rect 1086 152 1089 158
rect 1134 152 1137 168
rect 1054 142 1057 148
rect 930 128 934 131
rect 974 128 982 131
rect 942 111 945 118
rect 934 108 945 111
rect 934 82 937 108
rect 942 92 945 98
rect 950 72 953 108
rect 966 72 969 128
rect 906 58 913 61
rect 958 62 961 68
rect 870 52 873 58
rect 842 48 846 51
rect 722 28 726 31
rect 638 18 646 21
rect 622 -18 625 8
rect 646 -18 649 18
rect 694 -18 697 18
rect 782 -18 785 28
rect 806 -18 809 8
rect 838 -18 841 48
rect 878 11 881 58
rect 878 8 886 11
rect 886 -18 889 8
rect 902 -18 905 58
rect 974 12 977 128
rect 992 103 994 107
rect 998 103 1001 107
rect 1005 103 1008 107
rect 982 52 985 98
rect 994 78 998 81
rect 1022 62 1025 98
rect 1038 72 1041 78
rect 1030 62 1033 68
rect 1022 52 1025 58
rect 1054 52 1057 78
rect 982 -18 985 48
rect 1062 32 1065 148
rect 1102 102 1105 148
rect 1110 142 1113 148
rect 1150 122 1153 148
rect 1158 142 1161 148
rect 1182 142 1185 148
rect 1190 142 1193 218
rect 1198 181 1201 208
rect 1206 192 1209 258
rect 1230 212 1233 258
rect 1246 252 1249 258
rect 1198 178 1206 181
rect 1214 162 1217 168
rect 1190 122 1193 138
rect 1214 132 1217 138
rect 1046 -18 1049 8
rect 1070 -18 1073 78
rect 1110 72 1113 108
rect 1158 92 1161 98
rect 1126 72 1129 88
rect 1174 72 1177 118
rect 1214 82 1217 128
rect 1210 78 1214 81
rect 1182 72 1185 78
rect 1222 72 1225 168
rect 1246 142 1249 148
rect 1254 142 1257 298
rect 1262 262 1265 318
rect 1270 272 1273 278
rect 1282 268 1286 271
rect 1270 252 1273 258
rect 1290 248 1294 251
rect 1262 152 1265 238
rect 1286 152 1289 228
rect 1302 152 1305 258
rect 1310 201 1313 348
rect 1334 312 1337 348
rect 1366 312 1369 348
rect 1374 332 1377 338
rect 1350 292 1353 308
rect 1370 288 1374 291
rect 1318 262 1321 278
rect 1326 272 1329 288
rect 1382 282 1385 318
rect 1390 292 1393 348
rect 1406 342 1409 358
rect 1370 278 1374 281
rect 1338 268 1342 271
rect 1398 262 1401 338
rect 1414 281 1417 318
rect 1422 292 1425 318
rect 1430 282 1433 308
rect 1438 282 1441 368
rect 1446 362 1449 408
rect 1446 342 1449 358
rect 1462 342 1465 418
rect 1478 401 1481 458
rect 1486 442 1489 468
rect 1486 422 1489 438
rect 1478 398 1489 401
rect 1474 388 1478 391
rect 1486 352 1489 398
rect 1414 278 1425 281
rect 1322 258 1326 261
rect 1318 212 1321 218
rect 1310 198 1321 201
rect 1318 192 1321 198
rect 1350 182 1353 238
rect 1334 152 1337 158
rect 1342 152 1345 158
rect 1298 148 1302 151
rect 1354 148 1358 151
rect 1262 142 1265 148
rect 1286 142 1289 148
rect 1234 128 1238 131
rect 1238 92 1241 118
rect 1090 68 1094 71
rect 1242 68 1246 71
rect 1078 62 1081 68
rect 1090 58 1094 61
rect 1082 38 1086 41
rect 1102 32 1105 68
rect 1218 58 1222 61
rect 1250 58 1254 61
rect 1118 52 1121 58
rect 1234 48 1238 51
rect 1250 48 1254 51
rect 1262 51 1265 118
rect 1310 112 1313 148
rect 1290 78 1294 81
rect 1342 72 1345 138
rect 1358 132 1361 138
rect 1350 72 1353 78
rect 1366 72 1369 158
rect 1398 152 1401 258
rect 1406 252 1409 258
rect 1414 202 1417 268
rect 1422 262 1425 278
rect 1446 232 1449 338
rect 1458 328 1462 331
rect 1454 282 1457 318
rect 1470 312 1473 338
rect 1478 272 1481 278
rect 1486 272 1489 348
rect 1494 332 1497 458
rect 1510 452 1513 468
rect 1534 462 1537 538
rect 1514 448 1518 451
rect 1512 403 1514 407
rect 1518 403 1521 407
rect 1525 403 1528 407
rect 1526 342 1529 348
rect 1518 312 1521 318
rect 1526 282 1529 328
rect 1458 268 1462 271
rect 1474 268 1478 271
rect 1482 258 1486 261
rect 1494 261 1497 278
rect 1490 258 1497 261
rect 1454 242 1457 258
rect 1406 142 1409 168
rect 1414 152 1417 198
rect 1430 192 1433 198
rect 1450 178 1454 181
rect 1450 148 1454 151
rect 1386 138 1390 141
rect 1434 138 1438 141
rect 1374 132 1377 138
rect 1394 128 1398 131
rect 1382 122 1385 128
rect 1382 72 1385 98
rect 1398 82 1401 118
rect 1446 82 1449 138
rect 1454 132 1457 148
rect 1462 92 1465 248
rect 1470 162 1473 258
rect 1526 222 1529 278
rect 1534 242 1537 458
rect 1542 412 1545 728
rect 1566 721 1569 738
rect 1558 718 1569 721
rect 1550 622 1553 678
rect 1550 602 1553 618
rect 1558 582 1561 718
rect 1566 692 1569 708
rect 1574 612 1577 678
rect 1582 661 1585 738
rect 1590 682 1593 688
rect 1582 658 1590 661
rect 1574 592 1577 598
rect 1550 552 1553 568
rect 1590 552 1593 658
rect 1598 632 1601 938
rect 1606 892 1609 938
rect 1606 861 1609 888
rect 1614 882 1617 898
rect 1622 892 1625 938
rect 1670 901 1673 918
rect 1670 898 1681 901
rect 1622 872 1625 878
rect 1646 872 1649 878
rect 1606 858 1614 861
rect 1638 841 1641 858
rect 1630 838 1641 841
rect 1630 832 1633 838
rect 1642 828 1646 831
rect 1606 762 1609 768
rect 1614 752 1617 828
rect 1654 812 1657 888
rect 1670 882 1673 888
rect 1678 882 1681 898
rect 1686 892 1689 928
rect 1694 872 1697 938
rect 1702 872 1705 878
rect 1666 858 1673 861
rect 1670 852 1673 858
rect 1678 852 1681 858
rect 1718 851 1721 918
rect 1730 858 1734 861
rect 1718 848 1726 851
rect 1662 841 1665 848
rect 1686 841 1689 848
rect 1662 838 1689 841
rect 1654 802 1657 808
rect 1630 762 1633 768
rect 1638 762 1641 788
rect 1654 742 1657 768
rect 1694 752 1697 788
rect 1614 722 1617 738
rect 1654 722 1657 738
rect 1662 732 1665 748
rect 1686 742 1689 748
rect 1670 732 1673 738
rect 1622 702 1625 718
rect 1646 702 1649 718
rect 1662 682 1665 728
rect 1702 691 1705 808
rect 1710 742 1713 818
rect 1718 812 1721 848
rect 1742 752 1745 948
rect 1758 921 1761 1018
rect 1782 992 1785 1068
rect 1790 1012 1793 1068
rect 1806 962 1809 1058
rect 1814 1032 1817 1068
rect 1854 1062 1857 1138
rect 1862 1138 1873 1141
rect 1878 1142 1881 1178
rect 1862 1122 1865 1138
rect 1754 918 1761 921
rect 1766 882 1769 948
rect 1782 892 1785 958
rect 1802 948 1806 951
rect 1790 942 1793 948
rect 1798 882 1801 948
rect 1810 938 1814 941
rect 1754 868 1758 871
rect 1806 871 1809 908
rect 1802 868 1809 871
rect 1822 862 1825 868
rect 1830 862 1833 948
rect 1850 940 1854 943
rect 1862 942 1865 1088
rect 1870 1012 1873 1128
rect 1878 1082 1881 1128
rect 1886 1092 1889 1218
rect 1918 1178 1926 1181
rect 1918 1172 1921 1178
rect 1906 1168 1910 1171
rect 1958 1162 1961 1188
rect 1990 1162 1993 1228
rect 1998 1202 2001 1258
rect 2006 1252 2009 1268
rect 2022 1242 2025 1268
rect 2038 1222 2041 1228
rect 2014 1211 2017 1218
rect 2046 1212 2049 1268
rect 2058 1238 2065 1241
rect 2006 1208 2017 1211
rect 2006 1162 2009 1208
rect 1966 1152 1969 1158
rect 1938 1148 1950 1151
rect 1910 1122 1913 1148
rect 1982 1142 1985 1148
rect 1990 1142 1993 1148
rect 1926 1138 1934 1141
rect 1926 1132 1929 1138
rect 1938 1128 1942 1131
rect 1934 1092 1937 1118
rect 1958 1102 1961 1138
rect 1886 1072 1889 1078
rect 1886 1052 1889 1058
rect 1878 1042 1881 1048
rect 1878 992 1881 1028
rect 1886 972 1889 1018
rect 1894 962 1897 1088
rect 1974 1082 1977 1138
rect 1982 1112 1985 1138
rect 1998 1132 2001 1158
rect 2014 1142 2017 1198
rect 2022 1192 2025 1208
rect 2062 1192 2065 1238
rect 2070 1202 2073 1258
rect 2078 1241 2081 1268
rect 2110 1262 2113 1268
rect 2118 1262 2121 1308
rect 2126 1272 2129 1298
rect 2142 1292 2145 1318
rect 2158 1272 2161 1348
rect 2166 1332 2169 1338
rect 2134 1262 2137 1268
rect 2162 1258 2177 1261
rect 2162 1248 2166 1251
rect 2150 1242 2153 1248
rect 2078 1238 2102 1241
rect 2134 1212 2137 1228
rect 2006 1132 2009 1138
rect 2022 1131 2025 1138
rect 2014 1128 2025 1131
rect 2014 1121 2017 1128
rect 2010 1118 2017 1121
rect 2038 1122 2041 1158
rect 2024 1103 2026 1107
rect 2030 1103 2033 1107
rect 2037 1103 2040 1107
rect 1998 1081 2001 1098
rect 2046 1092 2049 1188
rect 2054 1132 2057 1158
rect 2062 1092 2065 1178
rect 2078 1152 2081 1208
rect 2118 1142 2121 1188
rect 2126 1182 2129 1188
rect 2106 1138 2110 1141
rect 2070 1112 2073 1138
rect 2010 1088 2014 1091
rect 1998 1078 2017 1081
rect 1902 1072 1905 1078
rect 1910 1072 1913 1078
rect 1902 1002 1905 1038
rect 1910 1002 1913 1068
rect 1934 1058 1942 1061
rect 1918 1052 1921 1058
rect 1934 1012 1937 1058
rect 1942 992 1945 1038
rect 1950 1022 1953 1058
rect 1966 1052 1969 1078
rect 2014 1072 2017 1078
rect 2030 1078 2049 1081
rect 2058 1078 2062 1081
rect 2030 1072 2033 1078
rect 2046 1072 2049 1078
rect 1986 1068 1990 1071
rect 1974 1062 1977 1068
rect 1998 1062 2001 1068
rect 2038 1062 2041 1068
rect 1874 948 1878 951
rect 1970 948 1974 951
rect 1838 912 1841 918
rect 1886 912 1889 928
rect 1846 862 1849 888
rect 1894 871 1897 948
rect 1910 942 1913 948
rect 1918 922 1921 948
rect 1946 938 1958 941
rect 1890 868 1897 871
rect 1762 858 1766 861
rect 1750 802 1753 818
rect 1766 752 1769 838
rect 1774 752 1777 858
rect 1806 832 1809 858
rect 1834 848 1838 851
rect 1794 788 1798 791
rect 1834 788 1838 791
rect 1814 762 1817 768
rect 1846 761 1849 818
rect 1878 802 1881 858
rect 1846 758 1854 761
rect 1834 748 1838 751
rect 1734 742 1737 748
rect 1742 732 1745 748
rect 1750 732 1753 738
rect 1694 688 1705 691
rect 1714 728 1718 731
rect 1610 678 1614 681
rect 1610 658 1614 661
rect 1642 658 1646 661
rect 1630 651 1633 658
rect 1630 648 1641 651
rect 1658 648 1662 651
rect 1614 592 1617 628
rect 1626 618 1630 621
rect 1638 592 1641 648
rect 1598 552 1601 558
rect 1590 512 1593 548
rect 1598 542 1601 548
rect 1586 488 1590 491
rect 1550 482 1553 488
rect 1542 352 1545 408
rect 1550 342 1553 418
rect 1566 372 1569 478
rect 1606 472 1609 578
rect 1650 568 1654 571
rect 1614 512 1617 518
rect 1630 472 1633 558
rect 1658 548 1662 551
rect 1638 542 1641 548
rect 1670 522 1673 668
rect 1678 662 1681 688
rect 1694 672 1697 688
rect 1710 681 1713 728
rect 1730 718 1734 721
rect 1722 688 1726 691
rect 1702 678 1713 681
rect 1722 678 1726 681
rect 1686 652 1689 658
rect 1694 652 1697 668
rect 1702 662 1705 678
rect 1714 668 1718 671
rect 1738 668 1742 671
rect 1750 652 1753 658
rect 1734 642 1737 648
rect 1694 562 1697 628
rect 1710 592 1713 608
rect 1750 562 1753 568
rect 1694 552 1697 558
rect 1742 552 1745 558
rect 1758 552 1761 718
rect 1766 682 1769 728
rect 1774 692 1777 748
rect 1862 742 1865 748
rect 1878 742 1881 748
rect 1886 742 1889 848
rect 1894 742 1897 858
rect 1902 822 1905 918
rect 1926 911 1929 938
rect 1918 908 1929 911
rect 1934 922 1937 928
rect 1942 922 1945 928
rect 1982 922 1985 958
rect 1990 952 1993 1058
rect 1998 952 2001 1048
rect 2006 962 2009 998
rect 2062 992 2065 1048
rect 2070 1002 2073 1108
rect 2086 1072 2089 1088
rect 2094 1072 2097 1118
rect 2102 1112 2105 1128
rect 2118 1082 2121 1088
rect 2106 1068 2113 1071
rect 2090 1058 2094 1061
rect 2098 1058 2105 1061
rect 2078 1052 2081 1058
rect 2094 992 2097 1048
rect 2102 982 2105 1058
rect 2110 1052 2113 1068
rect 2118 1062 2121 1068
rect 2126 1062 2129 1108
rect 2134 1092 2137 1148
rect 2142 1142 2145 1178
rect 2134 1078 2142 1081
rect 2022 942 2025 948
rect 2046 942 2049 968
rect 2062 948 2070 951
rect 2054 942 2057 948
rect 2062 932 2065 948
rect 2086 942 2089 968
rect 2074 938 2078 941
rect 2094 932 2097 948
rect 1918 872 1921 908
rect 1934 862 1937 918
rect 1950 872 1953 888
rect 1958 872 1961 878
rect 1974 872 1977 878
rect 1982 862 1985 918
rect 2006 872 2009 888
rect 1954 858 1958 861
rect 1994 858 1998 861
rect 2014 852 2017 918
rect 2024 903 2026 907
rect 2030 903 2033 907
rect 2037 903 2040 907
rect 1930 848 1934 851
rect 1970 848 1974 851
rect 1982 842 1985 848
rect 2038 842 2041 858
rect 1910 802 1913 818
rect 1834 738 1838 741
rect 1822 702 1825 738
rect 1778 668 1782 671
rect 1790 662 1793 698
rect 1818 688 1822 691
rect 1822 602 1825 678
rect 1830 662 1833 708
rect 1862 692 1865 718
rect 1886 692 1889 738
rect 1846 682 1849 688
rect 1854 672 1857 688
rect 1874 678 1881 681
rect 1850 658 1854 661
rect 1870 642 1873 658
rect 1878 592 1881 678
rect 1902 672 1905 798
rect 1910 762 1913 788
rect 1934 752 1937 808
rect 1942 792 1945 818
rect 1910 662 1913 678
rect 1926 662 1929 738
rect 1934 732 1937 748
rect 1942 742 1945 758
rect 1950 751 1953 798
rect 1998 792 2001 818
rect 2014 762 2017 788
rect 2046 762 2049 908
rect 2054 872 2057 918
rect 2066 868 2070 871
rect 2086 862 2089 868
rect 2066 858 2070 861
rect 2054 852 2057 858
rect 2082 848 2086 851
rect 2094 812 2097 918
rect 2110 862 2113 958
rect 2118 942 2121 948
rect 2134 932 2137 1078
rect 2150 1062 2153 1228
rect 2158 1172 2161 1238
rect 2174 1231 2177 1258
rect 2166 1228 2177 1231
rect 2166 1172 2169 1228
rect 2158 1142 2161 1168
rect 2174 1162 2177 1218
rect 2182 1201 2185 1358
rect 2198 1342 2201 1368
rect 2206 1352 2209 1458
rect 2222 1362 2225 1388
rect 2238 1361 2241 1448
rect 2254 1442 2257 1448
rect 2234 1358 2241 1361
rect 2230 1352 2233 1358
rect 2194 1328 2198 1331
rect 2198 1292 2201 1308
rect 2190 1262 2193 1288
rect 2206 1281 2209 1298
rect 2214 1292 2217 1338
rect 2230 1321 2233 1338
rect 2226 1318 2233 1321
rect 2238 1311 2241 1318
rect 2222 1308 2241 1311
rect 2222 1302 2225 1308
rect 2246 1301 2249 1428
rect 2254 1392 2257 1408
rect 2270 1392 2273 1478
rect 2286 1472 2289 1478
rect 2278 1402 2281 1458
rect 2294 1442 2297 1538
rect 2318 1492 2321 1528
rect 2310 1482 2313 1488
rect 2302 1478 2310 1481
rect 2302 1361 2305 1478
rect 2322 1458 2326 1461
rect 2310 1402 2313 1458
rect 2334 1381 2337 1628
rect 2350 1592 2353 1668
rect 2358 1642 2361 1658
rect 2358 1542 2361 1638
rect 2374 1632 2377 1658
rect 2374 1552 2377 1558
rect 2326 1378 2337 1381
rect 2342 1382 2345 1418
rect 2350 1392 2353 1498
rect 2358 1491 2361 1518
rect 2366 1502 2369 1538
rect 2382 1511 2385 1558
rect 2390 1552 2393 1708
rect 2398 1692 2401 1718
rect 2406 1681 2409 1738
rect 2406 1678 2414 1681
rect 2398 1672 2401 1678
rect 2422 1671 2425 1828
rect 2430 1822 2433 1838
rect 2442 1818 2446 1821
rect 2494 1812 2497 1818
rect 2558 1812 2561 1828
rect 2536 1803 2538 1807
rect 2542 1803 2545 1807
rect 2549 1803 2552 1807
rect 2454 1762 2457 1798
rect 2498 1768 2502 1771
rect 2442 1748 2446 1751
rect 2430 1722 2433 1728
rect 2438 1692 2441 1738
rect 2454 1732 2457 1748
rect 2462 1712 2465 1718
rect 2462 1672 2465 1678
rect 2470 1672 2473 1738
rect 2510 1732 2513 1788
rect 2566 1782 2569 1838
rect 2582 1822 2585 1848
rect 2598 1832 2601 1918
rect 2606 1862 2609 1908
rect 2614 1902 2617 1948
rect 2638 1942 2641 1948
rect 2686 1942 2689 1998
rect 2806 1992 2809 2038
rect 2746 1988 2750 1991
rect 2710 1962 2713 1968
rect 2726 1942 2729 1958
rect 2662 1922 2665 1928
rect 2694 1892 2697 1918
rect 2654 1882 2657 1888
rect 2626 1878 2630 1881
rect 2666 1878 2670 1881
rect 2686 1872 2689 1878
rect 2650 1868 2654 1871
rect 2674 1868 2678 1871
rect 2622 1862 2625 1868
rect 2662 1862 2665 1868
rect 2694 1861 2697 1878
rect 2702 1872 2705 1928
rect 2742 1922 2745 1968
rect 2758 1962 2761 1988
rect 2814 1952 2817 2018
rect 2822 1952 2825 2148
rect 2846 2142 2849 2268
rect 2862 2252 2865 2258
rect 2862 2202 2865 2218
rect 2866 2148 2870 2151
rect 2854 2142 2857 2148
rect 2834 2138 2838 2141
rect 2830 2092 2833 2098
rect 2838 1992 2841 2118
rect 2846 2062 2849 2108
rect 2854 2082 2857 2138
rect 2862 2122 2865 2138
rect 2862 2032 2865 2118
rect 2870 2062 2873 2128
rect 2870 2032 2873 2058
rect 2878 2052 2881 2308
rect 2922 2288 2926 2291
rect 2910 2272 2913 2278
rect 2934 2262 2937 2298
rect 2942 2272 2945 2338
rect 2982 2302 2985 2348
rect 2998 2302 3001 2338
rect 3010 2328 3014 2331
rect 2998 2272 3001 2278
rect 3006 2272 3009 2328
rect 3030 2292 3033 2438
rect 3038 2342 3041 2348
rect 3054 2332 3057 2408
rect 3070 2362 3073 2418
rect 3050 2318 3054 2321
rect 3040 2303 3042 2307
rect 3046 2303 3049 2307
rect 3053 2303 3056 2307
rect 2902 2252 2905 2258
rect 2886 2242 2889 2248
rect 2902 2192 2905 2248
rect 2918 2212 2921 2248
rect 2934 2192 2937 2258
rect 2942 2191 2945 2268
rect 2950 2252 2953 2268
rect 3054 2262 3057 2268
rect 3062 2262 3065 2268
rect 2950 2202 2953 2248
rect 2970 2218 2974 2221
rect 2998 2212 3001 2258
rect 3034 2248 3038 2251
rect 3066 2248 3070 2251
rect 3078 2242 3081 2448
rect 3094 2412 3097 2518
rect 3102 2472 3105 2498
rect 3110 2482 3113 2518
rect 3118 2492 3121 2518
rect 3102 2402 3105 2458
rect 3094 2382 3097 2388
rect 3090 2348 3094 2351
rect 3110 2342 3113 2478
rect 3118 2472 3121 2478
rect 3126 2472 3129 2498
rect 3142 2492 3145 2518
rect 3158 2492 3161 2508
rect 3194 2488 3198 2491
rect 3166 2482 3169 2488
rect 3174 2462 3177 2468
rect 3146 2458 3150 2461
rect 3118 2452 3121 2458
rect 3138 2448 3142 2451
rect 3182 2432 3185 2468
rect 3202 2448 3206 2451
rect 3118 2392 3121 2428
rect 3142 2342 3145 2368
rect 3214 2362 3217 2718
rect 3222 2671 3225 2738
rect 3234 2728 3238 2731
rect 3246 2722 3249 2858
rect 3254 2782 3257 2858
rect 3254 2752 3257 2778
rect 3262 2762 3265 2768
rect 3270 2731 3273 2868
rect 3286 2842 3289 2868
rect 3294 2852 3297 2858
rect 3310 2852 3313 2928
rect 3334 2882 3337 2948
rect 3322 2878 3326 2881
rect 3322 2868 3326 2871
rect 3342 2862 3345 3048
rect 3358 2992 3361 3048
rect 3350 2922 3353 2928
rect 3366 2912 3369 3068
rect 3422 2942 3425 3068
rect 3374 2932 3377 2938
rect 3422 2932 3425 2938
rect 3374 2892 3377 2928
rect 3398 2892 3401 2908
rect 3430 2892 3433 2948
rect 3438 2902 3441 3058
rect 3350 2882 3353 2888
rect 3446 2882 3449 2888
rect 3378 2878 3382 2881
rect 3438 2872 3441 2878
rect 3354 2868 3358 2871
rect 3418 2868 3422 2871
rect 3330 2858 3334 2861
rect 3354 2858 3358 2861
rect 3418 2858 3425 2861
rect 3286 2812 3289 2838
rect 3318 2832 3321 2838
rect 3318 2818 3326 2821
rect 3318 2792 3321 2818
rect 3334 2792 3337 2848
rect 3350 2842 3353 2848
rect 3406 2802 3409 2858
rect 3282 2758 3286 2761
rect 3282 2748 3286 2751
rect 3298 2748 3302 2751
rect 3310 2742 3313 2748
rect 3278 2732 3281 2738
rect 3270 2728 3278 2731
rect 3290 2718 3294 2721
rect 3270 2692 3273 2718
rect 3318 2692 3321 2778
rect 3358 2742 3361 2758
rect 3326 2722 3329 2728
rect 3306 2688 3310 2691
rect 3282 2678 3286 2681
rect 3222 2668 3233 2671
rect 3222 2612 3225 2658
rect 3230 2652 3233 2668
rect 3266 2668 3270 2671
rect 3246 2662 3249 2668
rect 3238 2622 3241 2628
rect 3246 2611 3249 2658
rect 3286 2652 3289 2668
rect 3334 2662 3337 2668
rect 3342 2662 3345 2728
rect 3350 2702 3353 2740
rect 3382 2731 3385 2748
rect 3398 2742 3401 2758
rect 3422 2752 3425 2858
rect 3446 2852 3449 2858
rect 3430 2762 3433 2768
rect 3446 2752 3449 2808
rect 3454 2802 3457 3218
rect 3478 3202 3481 3218
rect 3462 3122 3465 3148
rect 3502 3142 3505 3158
rect 3486 2972 3489 3018
rect 3470 2952 3473 2968
rect 3482 2948 3486 2951
rect 3502 2932 3505 3138
rect 3510 3092 3513 3248
rect 3522 3148 3526 3151
rect 3534 3142 3537 3148
rect 3518 2982 3521 3018
rect 3518 2952 3521 2968
rect 3518 2932 3521 2948
rect 3478 2882 3481 2928
rect 3510 2882 3513 2918
rect 3526 2902 3529 3078
rect 3534 2952 3537 3058
rect 3542 2972 3545 3218
rect 3550 3092 3553 3328
rect 3558 3142 3561 3148
rect 3546 2948 3550 2951
rect 3534 2912 3537 2918
rect 3534 2882 3537 2888
rect 3490 2878 3494 2881
rect 3522 2878 3526 2881
rect 3474 2868 3478 2871
rect 3538 2868 3542 2871
rect 3494 2862 3497 2868
rect 3502 2862 3505 2868
rect 3526 2862 3529 2868
rect 3546 2858 3550 2861
rect 3470 2782 3473 2858
rect 3478 2792 3481 2818
rect 3502 2792 3505 2858
rect 3514 2848 3518 2851
rect 3534 2772 3537 2778
rect 3474 2768 3478 2771
rect 3486 2752 3489 2768
rect 3502 2752 3505 2768
rect 3406 2742 3409 2748
rect 3394 2738 3398 2741
rect 3382 2728 3393 2731
rect 3358 2692 3361 2718
rect 3366 2692 3369 2718
rect 3390 2692 3393 2728
rect 3370 2678 3374 2681
rect 3386 2678 3390 2681
rect 3406 2672 3409 2708
rect 3414 2672 3417 2748
rect 3510 2742 3513 2748
rect 3426 2738 3433 2741
rect 3430 2692 3433 2738
rect 3446 2738 3454 2741
rect 3446 2722 3449 2738
rect 3462 2732 3465 2738
rect 3482 2728 3486 2731
rect 3518 2722 3521 2740
rect 3526 2732 3529 2758
rect 3542 2752 3545 2758
rect 3558 2742 3561 2748
rect 3446 2692 3449 2718
rect 3422 2682 3425 2688
rect 3430 2682 3433 2688
rect 3478 2682 3481 2688
rect 3342 2632 3345 2658
rect 3238 2608 3249 2611
rect 3222 2562 3225 2608
rect 3238 2592 3241 2608
rect 3286 2592 3289 2628
rect 3246 2582 3249 2588
rect 3222 2472 3225 2558
rect 3334 2552 3337 2618
rect 3342 2562 3345 2578
rect 3350 2572 3353 2668
rect 3390 2652 3393 2658
rect 3406 2652 3409 2668
rect 3414 2652 3417 2658
rect 3374 2602 3377 2618
rect 3366 2562 3369 2568
rect 3346 2558 3353 2561
rect 3282 2548 3286 2551
rect 3262 2532 3265 2538
rect 3242 2528 3246 2531
rect 3230 2481 3233 2528
rect 3230 2478 3238 2481
rect 3258 2468 3262 2471
rect 3222 2462 3225 2468
rect 3230 2432 3233 2468
rect 3250 2458 3254 2461
rect 3270 2452 3273 2548
rect 3310 2522 3313 2528
rect 3286 2512 3289 2518
rect 3310 2502 3313 2518
rect 3290 2488 3294 2491
rect 3310 2472 3313 2498
rect 3318 2462 3321 2548
rect 3350 2542 3353 2558
rect 3390 2552 3393 2648
rect 3398 2572 3401 2618
rect 3438 2612 3441 2678
rect 3486 2672 3489 2708
rect 3494 2682 3497 2698
rect 3526 2678 3529 2728
rect 3494 2672 3497 2678
rect 3558 2672 3561 2688
rect 3450 2668 3454 2671
rect 3514 2638 3518 2641
rect 3406 2592 3409 2608
rect 3422 2542 3425 2558
rect 3438 2542 3441 2598
rect 3462 2582 3465 2618
rect 3554 2578 3558 2581
rect 3342 2492 3345 2528
rect 3334 2478 3337 2488
rect 3366 2472 3369 2518
rect 3374 2482 3377 2538
rect 3422 2522 3425 2538
rect 3470 2492 3473 2548
rect 3426 2478 3430 2481
rect 3382 2472 3385 2478
rect 3394 2468 3398 2471
rect 3410 2458 3414 2461
rect 3278 2432 3281 2448
rect 3302 2442 3305 2458
rect 3370 2448 3374 2451
rect 3246 2372 3249 2418
rect 3294 2362 3297 2368
rect 3150 2358 3158 2361
rect 3234 2358 3238 2361
rect 3098 2338 3102 2341
rect 3126 2332 3129 2338
rect 3134 2302 3137 2318
rect 3130 2268 3134 2271
rect 3118 2262 3121 2268
rect 3090 2248 3094 2251
rect 3102 2222 3105 2258
rect 3134 2252 3137 2258
rect 2942 2188 2953 2191
rect 2934 2162 2937 2168
rect 2922 2158 2926 2161
rect 2890 2148 2894 2151
rect 2898 2138 2902 2141
rect 2910 2132 2913 2158
rect 2942 2152 2945 2158
rect 2918 2132 2921 2148
rect 2934 2132 2937 2148
rect 2942 2091 2945 2138
rect 2938 2088 2945 2091
rect 2886 2072 2889 2078
rect 2894 2062 2897 2088
rect 2906 2078 2910 2081
rect 2906 2068 2910 2071
rect 2922 2068 2926 2071
rect 2934 2062 2937 2088
rect 2918 2052 2921 2058
rect 2878 2022 2881 2048
rect 2942 2042 2945 2048
rect 2950 2032 2953 2188
rect 2974 2182 2977 2188
rect 3106 2178 3110 2181
rect 2962 2158 2966 2161
rect 3010 2158 3014 2161
rect 2958 2132 2961 2138
rect 2966 2092 2969 2138
rect 2990 2132 2993 2158
rect 2998 2132 3001 2138
rect 2894 1992 2897 2028
rect 2958 2022 2961 2058
rect 2966 2032 2969 2068
rect 2974 2052 2977 2078
rect 3022 2062 3025 2178
rect 3142 2171 3145 2338
rect 3150 2292 3153 2358
rect 3162 2348 3166 2351
rect 3174 2342 3177 2358
rect 3254 2352 3257 2358
rect 3326 2352 3329 2358
rect 3186 2348 3190 2351
rect 3162 2338 3166 2341
rect 3202 2338 3206 2341
rect 3158 2272 3161 2278
rect 3158 2262 3161 2268
rect 3150 2242 3153 2248
rect 3166 2192 3169 2308
rect 3174 2302 3177 2338
rect 3174 2292 3177 2298
rect 3214 2292 3217 2348
rect 3238 2332 3241 2338
rect 3226 2328 3230 2331
rect 3246 2312 3249 2318
rect 3254 2312 3257 2348
rect 3334 2342 3337 2368
rect 3342 2352 3345 2448
rect 3390 2392 3393 2448
rect 3454 2422 3457 2458
rect 3470 2452 3473 2468
rect 3438 2362 3441 2368
rect 3402 2358 3406 2361
rect 3466 2358 3470 2361
rect 3314 2338 3318 2341
rect 3174 2222 3177 2248
rect 3182 2242 3185 2268
rect 3190 2262 3193 2268
rect 3182 2192 3185 2218
rect 3142 2168 3150 2171
rect 3070 2162 3073 2168
rect 3150 2162 3153 2168
rect 3166 2162 3169 2188
rect 3190 2182 3193 2218
rect 3198 2161 3201 2288
rect 3214 2272 3217 2278
rect 3262 2272 3265 2338
rect 3310 2322 3313 2338
rect 3350 2332 3353 2348
rect 3358 2342 3361 2358
rect 3382 2352 3385 2358
rect 3414 2342 3417 2348
rect 3386 2338 3390 2341
rect 3434 2338 3438 2341
rect 3322 2328 3326 2331
rect 3214 2252 3217 2258
rect 3206 2242 3209 2248
rect 3222 2242 3225 2248
rect 3238 2242 3241 2248
rect 3222 2212 3225 2238
rect 3246 2222 3249 2268
rect 3262 2222 3265 2248
rect 3270 2192 3273 2318
rect 3334 2312 3337 2328
rect 3334 2292 3337 2308
rect 3314 2288 3318 2291
rect 3358 2291 3361 2338
rect 3366 2332 3369 2338
rect 3378 2328 3382 2331
rect 3414 2322 3417 2338
rect 3422 2312 3425 2338
rect 3442 2328 3446 2331
rect 3454 2312 3457 2348
rect 3478 2342 3481 2348
rect 3390 2292 3393 2308
rect 3354 2288 3361 2291
rect 3350 2282 3353 2288
rect 3306 2268 3310 2271
rect 3286 2242 3289 2258
rect 3318 2242 3321 2248
rect 3342 2232 3345 2268
rect 3374 2262 3377 2288
rect 3398 2272 3401 2278
rect 3394 2248 3398 2251
rect 3390 2192 3393 2218
rect 3238 2162 3241 2168
rect 3198 2158 3206 2161
rect 3234 2158 3238 2161
rect 3290 2158 3294 2161
rect 3070 2142 3073 2148
rect 3086 2142 3089 2158
rect 3286 2152 3289 2158
rect 3154 2148 3158 2151
rect 3194 2148 3198 2151
rect 3218 2148 3222 2151
rect 3246 2148 3254 2151
rect 3030 2122 3033 2138
rect 3040 2103 3042 2107
rect 3046 2103 3049 2107
rect 3053 2103 3056 2107
rect 3034 2068 3038 2071
rect 3046 2062 3049 2078
rect 3054 2072 3057 2088
rect 3070 2082 3073 2138
rect 3078 2122 3081 2138
rect 3134 2132 3137 2138
rect 3078 2092 3081 2118
rect 3082 2078 3086 2081
rect 3070 2072 3073 2078
rect 3102 2072 3105 2078
rect 2986 2048 2990 2051
rect 2998 2042 3001 2058
rect 3054 2052 3057 2068
rect 3006 2042 3009 2048
rect 2942 1992 2945 2018
rect 2862 1962 2865 1988
rect 2846 1952 2849 1958
rect 2770 1948 2774 1951
rect 2750 1922 2753 1948
rect 2770 1938 2774 1941
rect 2710 1882 2713 1918
rect 2718 1871 2721 1888
rect 2714 1868 2721 1871
rect 2694 1858 2702 1861
rect 2738 1858 2742 1861
rect 2610 1838 2617 1841
rect 2598 1802 2601 1818
rect 2538 1748 2542 1751
rect 2574 1732 2577 1748
rect 2598 1742 2601 1748
rect 2590 1732 2593 1738
rect 2414 1668 2425 1671
rect 2402 1648 2406 1651
rect 2414 1562 2417 1668
rect 2422 1612 2425 1658
rect 2430 1621 2433 1668
rect 2438 1632 2441 1648
rect 2454 1632 2457 1668
rect 2486 1662 2489 1698
rect 2502 1672 2505 1708
rect 2494 1662 2497 1668
rect 2510 1662 2513 1718
rect 2558 1712 2561 1718
rect 2542 1682 2545 1698
rect 2474 1658 2478 1661
rect 2522 1658 2526 1661
rect 2542 1652 2545 1678
rect 2550 1672 2553 1688
rect 2554 1658 2558 1661
rect 2566 1651 2569 1728
rect 2574 1692 2577 1698
rect 2582 1692 2585 1718
rect 2598 1702 2601 1738
rect 2594 1678 2598 1681
rect 2582 1672 2585 1678
rect 2606 1662 2609 1718
rect 2614 1692 2617 1838
rect 2622 1722 2625 1848
rect 2638 1812 2641 1858
rect 2622 1672 2625 1678
rect 2630 1672 2633 1808
rect 2654 1792 2657 1798
rect 2662 1771 2665 1858
rect 2670 1791 2673 1818
rect 2678 1802 2681 1858
rect 2710 1851 2713 1858
rect 2702 1848 2713 1851
rect 2738 1848 2742 1851
rect 2702 1842 2705 1848
rect 2710 1832 2713 1848
rect 2750 1832 2753 1868
rect 2758 1852 2761 1858
rect 2670 1788 2678 1791
rect 2654 1768 2665 1771
rect 2654 1752 2657 1768
rect 2662 1752 2665 1758
rect 2642 1728 2646 1731
rect 2670 1692 2673 1778
rect 2678 1712 2681 1748
rect 2686 1712 2689 1738
rect 2694 1732 2697 1738
rect 2678 1672 2681 1678
rect 2686 1672 2689 1678
rect 2574 1658 2582 1661
rect 2654 1652 2657 1658
rect 2558 1648 2569 1651
rect 2430 1618 2441 1621
rect 2438 1592 2441 1618
rect 2454 1592 2457 1628
rect 2422 1572 2425 1588
rect 2374 1508 2385 1511
rect 2374 1491 2377 1508
rect 2358 1488 2377 1491
rect 2398 1492 2401 1548
rect 2414 1542 2417 1548
rect 2430 1542 2433 1588
rect 2422 1538 2430 1541
rect 2406 1532 2409 1538
rect 2422 1531 2425 1538
rect 2414 1528 2425 1531
rect 2446 1532 2449 1538
rect 2454 1532 2457 1548
rect 2462 1542 2465 1648
rect 2558 1632 2561 1648
rect 2574 1642 2577 1648
rect 2606 1642 2609 1648
rect 2638 1642 2641 1648
rect 2486 1612 2489 1618
rect 2536 1603 2538 1607
rect 2542 1603 2545 1607
rect 2549 1603 2552 1607
rect 2490 1588 2494 1591
rect 2482 1568 2494 1571
rect 2546 1568 2550 1571
rect 2510 1562 2513 1568
rect 2558 1562 2561 1628
rect 2358 1462 2361 1478
rect 2366 1402 2369 1478
rect 2302 1358 2313 1361
rect 2254 1332 2257 1348
rect 2262 1342 2265 1348
rect 2238 1298 2249 1301
rect 2238 1292 2241 1298
rect 2262 1292 2265 1298
rect 2206 1278 2217 1281
rect 2214 1272 2217 1278
rect 2242 1268 2246 1271
rect 2206 1262 2209 1268
rect 2190 1232 2193 1248
rect 2206 1202 2209 1258
rect 2262 1252 2265 1278
rect 2270 1262 2273 1348
rect 2294 1332 2297 1348
rect 2294 1292 2297 1328
rect 2302 1292 2305 1328
rect 2290 1278 2294 1281
rect 2310 1281 2313 1358
rect 2326 1352 2329 1378
rect 2342 1371 2345 1378
rect 2334 1368 2345 1371
rect 2374 1372 2377 1418
rect 2318 1312 2321 1348
rect 2334 1332 2337 1368
rect 2342 1352 2345 1358
rect 2358 1352 2361 1358
rect 2302 1278 2313 1281
rect 2342 1281 2345 1318
rect 2366 1312 2369 1338
rect 2382 1332 2385 1398
rect 2390 1352 2393 1478
rect 2406 1472 2409 1478
rect 2414 1462 2417 1528
rect 2446 1522 2449 1528
rect 2454 1472 2457 1518
rect 2434 1468 2438 1471
rect 2446 1468 2454 1471
rect 2422 1462 2425 1468
rect 2410 1458 2414 1461
rect 2430 1452 2433 1458
rect 2414 1412 2417 1448
rect 2414 1392 2417 1408
rect 2426 1348 2430 1351
rect 2406 1342 2409 1348
rect 2378 1328 2382 1331
rect 2374 1292 2377 1308
rect 2382 1292 2385 1318
rect 2390 1302 2393 1338
rect 2446 1332 2449 1468
rect 2454 1452 2457 1458
rect 2462 1452 2465 1478
rect 2470 1442 2473 1448
rect 2478 1362 2481 1478
rect 2486 1472 2489 1508
rect 2430 1292 2433 1298
rect 2406 1282 2409 1288
rect 2438 1282 2441 1288
rect 2462 1282 2465 1288
rect 2470 1282 2473 1328
rect 2478 1312 2481 1348
rect 2486 1322 2489 1458
rect 2502 1392 2505 1548
rect 2526 1532 2529 1538
rect 2518 1522 2521 1528
rect 2534 1492 2537 1498
rect 2550 1471 2553 1558
rect 2570 1548 2574 1551
rect 2558 1542 2561 1548
rect 2598 1542 2601 1548
rect 2606 1542 2609 1568
rect 2630 1552 2633 1578
rect 2654 1552 2657 1558
rect 2662 1552 2665 1648
rect 2678 1642 2681 1668
rect 2694 1612 2697 1658
rect 2678 1542 2681 1588
rect 2686 1542 2689 1548
rect 2582 1532 2585 1538
rect 2594 1528 2598 1531
rect 2642 1528 2646 1531
rect 2650 1528 2657 1531
rect 2558 1482 2561 1498
rect 2582 1492 2585 1498
rect 2590 1482 2593 1498
rect 2550 1468 2558 1471
rect 2514 1458 2518 1461
rect 2510 1412 2513 1448
rect 2558 1442 2561 1458
rect 2536 1403 2538 1407
rect 2542 1403 2545 1407
rect 2549 1403 2552 1407
rect 2510 1392 2513 1398
rect 2498 1358 2502 1361
rect 2510 1352 2513 1368
rect 2526 1351 2529 1368
rect 2546 1358 2550 1361
rect 2522 1348 2529 1351
rect 2498 1328 2502 1331
rect 2342 1278 2350 1281
rect 2494 1281 2497 1328
rect 2514 1288 2518 1291
rect 2534 1282 2537 1318
rect 2558 1292 2561 1408
rect 2582 1352 2585 1478
rect 2598 1462 2601 1468
rect 2606 1462 2609 1468
rect 2614 1392 2617 1518
rect 2622 1492 2625 1528
rect 2638 1502 2641 1518
rect 2630 1462 2633 1488
rect 2622 1362 2625 1368
rect 2602 1358 2606 1361
rect 2614 1352 2617 1358
rect 2570 1348 2574 1351
rect 2566 1332 2569 1348
rect 2638 1342 2641 1398
rect 2654 1352 2657 1528
rect 2662 1522 2665 1538
rect 2670 1522 2673 1528
rect 2678 1502 2681 1528
rect 2686 1482 2689 1488
rect 2670 1471 2673 1478
rect 2670 1468 2678 1471
rect 2662 1462 2665 1468
rect 2678 1462 2681 1468
rect 2666 1448 2670 1451
rect 2682 1448 2686 1451
rect 2574 1332 2577 1338
rect 2582 1332 2585 1338
rect 2582 1282 2585 1308
rect 2490 1278 2497 1281
rect 2522 1278 2526 1281
rect 2286 1252 2289 1258
rect 2230 1222 2233 1248
rect 2182 1198 2193 1201
rect 2190 1152 2193 1198
rect 2214 1192 2217 1198
rect 2230 1152 2233 1218
rect 2238 1192 2241 1248
rect 2294 1232 2297 1268
rect 2270 1152 2273 1218
rect 2274 1148 2278 1151
rect 2174 1142 2177 1148
rect 2198 1142 2201 1148
rect 2158 1062 2161 1068
rect 2142 1002 2145 1058
rect 2142 952 2145 998
rect 2150 942 2153 1058
rect 2166 1042 2169 1138
rect 2182 1092 2185 1138
rect 2206 1132 2209 1148
rect 2214 1142 2217 1148
rect 2262 1142 2265 1148
rect 2250 1138 2254 1141
rect 2230 1082 2233 1138
rect 2178 1078 2182 1081
rect 2238 1072 2241 1128
rect 2246 1082 2249 1098
rect 2262 1072 2265 1138
rect 2210 1068 2214 1071
rect 2174 1042 2177 1048
rect 2182 972 2185 1048
rect 2230 1042 2233 1058
rect 2182 958 2190 961
rect 2182 952 2185 958
rect 2198 952 2201 1018
rect 2250 988 2254 991
rect 2222 952 2225 968
rect 2230 952 2233 968
rect 2162 948 2166 951
rect 2262 942 2265 1068
rect 2278 1052 2281 1138
rect 2294 1092 2297 1228
rect 2302 1222 2305 1278
rect 2310 1211 2313 1268
rect 2318 1262 2321 1278
rect 2326 1252 2329 1258
rect 2326 1232 2329 1248
rect 2302 1208 2313 1211
rect 2302 1082 2305 1208
rect 2314 1158 2318 1161
rect 2318 1122 2321 1128
rect 2286 1062 2289 1068
rect 2310 1062 2313 1098
rect 2326 1082 2329 1218
rect 2334 1172 2337 1268
rect 2382 1262 2385 1278
rect 2342 1248 2350 1251
rect 2342 1192 2345 1248
rect 2374 1182 2377 1248
rect 2370 1148 2374 1151
rect 2350 1102 2353 1128
rect 2366 1122 2369 1138
rect 2350 1072 2353 1088
rect 2318 1068 2337 1071
rect 2318 1062 2321 1068
rect 2334 1062 2337 1068
rect 2358 1062 2361 1118
rect 2382 1082 2385 1148
rect 2310 1052 2313 1058
rect 2326 1052 2329 1058
rect 2290 1048 2294 1051
rect 2178 938 2182 941
rect 2134 892 2137 928
rect 2150 902 2153 918
rect 2122 868 2126 871
rect 2142 868 2150 871
rect 2162 868 2166 871
rect 2174 870 2177 898
rect 2182 871 2185 928
rect 2198 902 2201 928
rect 2194 888 2198 891
rect 2106 858 2110 861
rect 2114 858 2121 861
rect 2110 842 2113 848
rect 2066 768 2081 771
rect 1998 758 2006 761
rect 2078 761 2081 768
rect 2078 758 2094 761
rect 1990 752 1993 758
rect 1950 748 1961 751
rect 1958 742 1961 748
rect 1946 738 1950 741
rect 1986 738 1990 741
rect 1954 728 1958 731
rect 1974 722 1977 728
rect 1998 722 2001 758
rect 2030 742 2033 748
rect 2070 742 2073 758
rect 2082 748 2086 751
rect 2010 728 2014 731
rect 2098 728 2102 731
rect 2054 722 2057 728
rect 2062 722 2065 728
rect 1942 692 1945 708
rect 1950 672 1953 678
rect 2006 672 2009 678
rect 2014 672 2017 718
rect 2102 712 2105 718
rect 2024 703 2026 707
rect 2030 703 2033 707
rect 2037 703 2040 707
rect 2110 692 2113 808
rect 2118 752 2121 858
rect 2126 852 2129 858
rect 2134 842 2137 868
rect 2142 862 2145 868
rect 2182 868 2198 871
rect 2206 862 2209 868
rect 2222 862 2225 938
rect 2238 881 2241 928
rect 2234 878 2241 881
rect 2230 872 2233 878
rect 2154 858 2158 861
rect 2214 858 2222 861
rect 2150 802 2153 818
rect 2158 771 2161 858
rect 2206 792 2209 818
rect 2158 768 2169 771
rect 2166 762 2169 768
rect 2154 758 2158 761
rect 2130 748 2134 751
rect 2126 732 2129 738
rect 2134 722 2137 738
rect 2078 672 2081 678
rect 2026 668 2030 671
rect 1958 661 1961 668
rect 1950 658 1961 661
rect 2050 658 2054 661
rect 2074 658 2078 661
rect 1922 638 1926 641
rect 1934 641 1937 648
rect 1934 638 1942 641
rect 1886 572 1889 638
rect 1778 558 1782 561
rect 1798 552 1801 568
rect 1810 558 1814 561
rect 1770 548 1774 551
rect 1686 542 1689 548
rect 1714 538 1718 541
rect 1686 532 1689 538
rect 1710 522 1713 528
rect 1678 482 1681 488
rect 1578 468 1582 471
rect 1598 462 1601 468
rect 1614 462 1617 468
rect 1646 462 1649 468
rect 1582 442 1585 448
rect 1622 422 1625 458
rect 1638 452 1641 458
rect 1638 392 1641 418
rect 1610 348 1614 351
rect 1542 302 1545 338
rect 1582 312 1585 318
rect 1598 282 1601 338
rect 1610 328 1614 331
rect 1610 278 1614 281
rect 1550 272 1553 278
rect 1582 272 1585 278
rect 1570 268 1574 271
rect 1542 262 1545 268
rect 1550 251 1553 258
rect 1542 248 1553 251
rect 1570 248 1574 251
rect 1542 242 1545 248
rect 1582 222 1585 268
rect 1606 262 1609 268
rect 1598 252 1601 258
rect 1482 148 1486 151
rect 1502 151 1505 218
rect 1512 203 1514 207
rect 1518 203 1521 207
rect 1525 203 1528 207
rect 1534 152 1537 218
rect 1590 162 1593 218
rect 1606 192 1609 238
rect 1622 232 1625 348
rect 1630 342 1633 378
rect 1646 362 1649 458
rect 1654 422 1657 468
rect 1662 452 1665 458
rect 1670 442 1673 478
rect 1686 452 1689 458
rect 1694 422 1697 468
rect 1710 462 1713 468
rect 1678 372 1681 378
rect 1646 282 1649 358
rect 1662 312 1665 358
rect 1670 351 1673 368
rect 1670 348 1678 351
rect 1646 272 1649 278
rect 1646 262 1649 268
rect 1670 262 1673 318
rect 1678 272 1681 348
rect 1686 322 1689 338
rect 1694 332 1697 348
rect 1710 342 1713 458
rect 1718 392 1721 458
rect 1726 402 1729 548
rect 1798 522 1801 538
rect 1754 488 1758 491
rect 1778 458 1782 461
rect 1758 452 1761 458
rect 1790 452 1793 508
rect 1806 471 1809 558
rect 1822 502 1825 548
rect 1830 492 1833 538
rect 1838 492 1841 558
rect 1846 472 1849 538
rect 1862 532 1865 568
rect 1870 552 1873 558
rect 1878 522 1881 548
rect 1858 518 1862 521
rect 1894 502 1897 618
rect 1918 552 1921 558
rect 1926 552 1929 558
rect 1902 542 1905 548
rect 1910 542 1913 548
rect 1934 542 1937 598
rect 1950 562 1953 658
rect 2014 652 2017 658
rect 2050 648 2054 651
rect 2070 642 2073 648
rect 2086 642 2089 668
rect 2130 658 2134 661
rect 2094 652 2097 658
rect 2142 652 2145 758
rect 2166 752 2169 758
rect 2194 748 2198 751
rect 2158 692 2161 748
rect 2166 692 2169 748
rect 2214 742 2217 858
rect 2226 848 2230 851
rect 2254 812 2257 848
rect 2262 842 2265 918
rect 2270 892 2273 998
rect 2278 952 2281 1008
rect 2302 992 2305 1038
rect 2274 868 2278 871
rect 2286 862 2289 978
rect 2294 882 2297 918
rect 2302 912 2305 918
rect 2310 882 2313 1038
rect 2334 972 2337 1018
rect 2358 972 2361 1018
rect 2366 962 2369 1078
rect 2378 1058 2382 1061
rect 2390 992 2393 1268
rect 2422 1262 2425 1268
rect 2442 1258 2446 1261
rect 2466 1258 2470 1261
rect 2406 1162 2409 1218
rect 2414 1192 2417 1258
rect 2478 1252 2481 1258
rect 2486 1242 2489 1278
rect 2498 1268 2502 1271
rect 2494 1222 2497 1258
rect 2430 1182 2433 1218
rect 2446 1212 2449 1218
rect 2526 1202 2529 1268
rect 2542 1252 2545 1268
rect 2550 1252 2553 1258
rect 2536 1203 2538 1207
rect 2542 1203 2545 1207
rect 2549 1203 2552 1207
rect 2558 1192 2561 1238
rect 2414 1152 2417 1158
rect 2446 1142 2449 1178
rect 2402 1138 2406 1141
rect 2502 1142 2505 1168
rect 2510 1142 2513 1148
rect 2518 1142 2521 1148
rect 2454 1132 2457 1140
rect 2486 1132 2489 1138
rect 2526 1132 2529 1138
rect 2546 1128 2550 1131
rect 2478 1118 2486 1121
rect 2430 1092 2433 1118
rect 2398 1052 2401 1078
rect 2430 1062 2433 1068
rect 2478 1062 2481 1118
rect 2418 1058 2422 1061
rect 2406 1012 2409 1048
rect 2382 952 2385 958
rect 2330 948 2334 951
rect 2338 938 2342 941
rect 2374 942 2377 948
rect 2306 878 2310 881
rect 2318 881 2321 918
rect 2318 878 2329 881
rect 2314 868 2318 871
rect 2326 862 2329 878
rect 2342 862 2345 898
rect 2350 891 2353 918
rect 2366 912 2369 940
rect 2410 938 2414 941
rect 2350 888 2361 891
rect 2350 872 2353 878
rect 2358 862 2361 888
rect 2294 852 2297 858
rect 2342 852 2345 858
rect 2326 842 2329 848
rect 2222 752 2225 758
rect 2262 751 2265 838
rect 2258 748 2265 751
rect 2282 748 2286 751
rect 2246 742 2249 748
rect 2294 742 2297 758
rect 2342 751 2345 758
rect 2310 742 2313 748
rect 2226 738 2230 741
rect 2282 738 2286 741
rect 2174 722 2177 738
rect 2214 732 2217 738
rect 2250 728 2257 731
rect 2182 682 2185 718
rect 2254 701 2257 728
rect 2262 712 2265 738
rect 2278 722 2281 728
rect 2310 712 2313 728
rect 2254 698 2265 701
rect 2210 678 2214 681
rect 2150 662 2153 668
rect 2166 642 2169 678
rect 2186 668 2190 671
rect 2130 638 2134 641
rect 2174 622 2177 658
rect 2198 652 2201 658
rect 1982 562 1985 598
rect 1990 581 1993 618
rect 2110 582 2113 598
rect 1990 578 1998 581
rect 2110 562 2113 578
rect 1994 558 1998 561
rect 2010 558 2017 561
rect 1950 542 1953 558
rect 1962 538 1966 541
rect 1910 531 1913 538
rect 1982 531 1985 558
rect 2014 552 2017 558
rect 2074 558 2078 561
rect 2122 558 2126 561
rect 2046 552 2049 558
rect 2002 548 2006 551
rect 1902 528 1913 531
rect 1974 528 1985 531
rect 1874 478 1878 481
rect 1802 468 1809 471
rect 1734 392 1737 448
rect 1778 438 1782 441
rect 1718 352 1721 388
rect 1742 352 1745 438
rect 1806 432 1809 458
rect 1818 448 1822 451
rect 1750 352 1753 368
rect 1738 348 1742 351
rect 1710 332 1713 338
rect 1702 301 1705 318
rect 1726 312 1729 328
rect 1702 298 1713 301
rect 1698 288 1702 291
rect 1710 291 1713 298
rect 1750 292 1753 338
rect 1710 288 1721 291
rect 1702 278 1710 281
rect 1686 272 1689 278
rect 1718 271 1721 288
rect 1758 282 1761 348
rect 1766 331 1769 418
rect 1774 392 1777 398
rect 1822 392 1825 438
rect 1778 348 1782 351
rect 1790 342 1793 358
rect 1810 348 1814 351
rect 1822 342 1825 348
rect 1766 328 1774 331
rect 1798 328 1806 331
rect 1790 292 1793 318
rect 1762 278 1766 281
rect 1718 268 1726 271
rect 1742 262 1745 268
rect 1766 262 1769 268
rect 1798 262 1801 318
rect 1814 292 1817 308
rect 1830 292 1833 468
rect 1846 442 1849 468
rect 1846 362 1849 438
rect 1854 392 1857 458
rect 1846 352 1849 358
rect 1854 352 1857 388
rect 1838 342 1841 348
rect 1862 341 1865 458
rect 1854 338 1865 341
rect 1634 258 1638 261
rect 1722 258 1726 261
rect 1650 248 1654 251
rect 1674 248 1678 251
rect 1630 192 1633 248
rect 1638 162 1641 218
rect 1554 158 1558 161
rect 1542 152 1545 158
rect 1502 148 1513 151
rect 1590 148 1606 151
rect 1498 138 1502 141
rect 1486 122 1489 138
rect 1510 132 1513 148
rect 1526 132 1529 138
rect 1498 78 1502 81
rect 1290 68 1294 71
rect 1274 58 1278 61
rect 1322 58 1326 61
rect 1262 48 1270 51
rect 1214 -18 1217 8
rect 1270 -18 1273 8
rect 518 -19 522 -18
rect 510 -22 522 -19
rect 606 -22 610 -18
rect 622 -22 626 -18
rect 646 -22 650 -18
rect 694 -22 698 -18
rect 782 -22 786 -18
rect 806 -22 810 -18
rect 838 -22 842 -18
rect 886 -22 890 -18
rect 902 -22 906 -18
rect 982 -22 986 -18
rect 1046 -22 1050 -18
rect 1070 -22 1074 -18
rect 1214 -22 1218 -18
rect 1270 -22 1274 -18
rect 1334 -19 1338 -18
rect 1342 -19 1345 68
rect 1354 58 1358 61
rect 1374 52 1377 58
rect 1398 52 1401 78
rect 1406 52 1409 68
rect 1414 62 1417 78
rect 1434 68 1438 71
rect 1426 58 1430 61
rect 1442 58 1446 61
rect 1462 52 1465 78
rect 1486 72 1489 78
rect 1514 68 1518 71
rect 1470 62 1473 68
rect 1478 62 1481 68
rect 1534 62 1537 98
rect 1542 72 1545 148
rect 1550 122 1553 148
rect 1590 142 1593 148
rect 1562 138 1566 141
rect 1586 128 1590 131
rect 1558 82 1561 128
rect 1598 92 1601 138
rect 1614 122 1617 138
rect 1638 102 1641 128
rect 1614 72 1617 78
rect 1522 58 1526 61
rect 1434 48 1438 51
rect 1566 42 1569 68
rect 1562 18 1566 21
rect 1614 12 1617 68
rect 1622 52 1625 58
rect 1638 52 1641 78
rect 1646 22 1649 158
rect 1654 142 1657 238
rect 1662 192 1665 228
rect 1678 192 1681 218
rect 1666 148 1670 151
rect 1654 72 1657 138
rect 1662 92 1665 138
rect 1670 102 1673 138
rect 1678 132 1681 158
rect 1702 152 1705 258
rect 1726 152 1729 198
rect 1694 142 1697 148
rect 1706 128 1710 131
rect 1726 92 1729 118
rect 1734 102 1737 258
rect 1774 252 1777 258
rect 1790 192 1793 258
rect 1806 252 1809 268
rect 1822 252 1825 278
rect 1830 192 1833 248
rect 1838 202 1841 308
rect 1854 302 1857 338
rect 1870 332 1873 428
rect 1878 382 1881 448
rect 1878 342 1881 378
rect 1886 332 1889 478
rect 1894 472 1897 478
rect 1902 452 1905 528
rect 1914 458 1918 461
rect 1910 442 1913 448
rect 1918 432 1921 458
rect 1926 452 1929 518
rect 1934 472 1937 498
rect 1950 471 1953 518
rect 1974 512 1977 528
rect 1986 518 1990 521
rect 1982 472 1985 498
rect 1998 472 2001 538
rect 2006 492 2009 538
rect 2014 492 2017 538
rect 2062 532 2065 538
rect 2090 528 2094 531
rect 2054 522 2057 528
rect 2024 503 2026 507
rect 2030 503 2033 507
rect 2037 503 2040 507
rect 2102 492 2105 528
rect 2050 478 2054 481
rect 1950 468 1961 471
rect 1950 452 1953 458
rect 1958 452 1961 468
rect 2002 468 2006 471
rect 1970 458 1974 461
rect 1918 402 1921 418
rect 1894 362 1897 378
rect 1894 352 1897 358
rect 1902 352 1905 368
rect 1926 342 1929 408
rect 1942 382 1945 418
rect 1950 372 1953 448
rect 1974 442 1977 448
rect 1982 371 1985 468
rect 1990 462 1993 468
rect 2014 392 2017 468
rect 2022 462 2025 468
rect 2022 422 2025 458
rect 1982 368 1993 371
rect 1990 362 1993 368
rect 2006 362 2009 378
rect 1946 358 1950 361
rect 1974 352 1977 358
rect 1982 352 1985 358
rect 2030 352 2033 478
rect 2062 471 2065 478
rect 2058 468 2065 471
rect 2086 472 2089 478
rect 2066 458 2070 461
rect 2054 452 2057 458
rect 2078 452 2081 458
rect 2026 348 2030 351
rect 1950 342 1953 348
rect 2006 342 2009 348
rect 1914 328 1918 331
rect 1862 312 1865 318
rect 1854 272 1857 288
rect 1862 282 1865 288
rect 1862 272 1865 278
rect 1846 242 1849 258
rect 1870 252 1873 258
rect 1878 242 1881 268
rect 1886 262 1889 268
rect 1894 261 1897 318
rect 1910 312 1913 318
rect 1942 311 1945 318
rect 1942 308 1953 311
rect 1902 272 1905 298
rect 1942 292 1945 298
rect 1950 272 1953 308
rect 1966 282 1969 338
rect 1998 332 2001 338
rect 2022 332 2025 338
rect 2046 322 2049 358
rect 1914 268 1918 271
rect 1942 268 1950 271
rect 1894 258 1905 261
rect 1902 252 1905 258
rect 1890 248 1894 251
rect 1910 242 1913 258
rect 1926 252 1929 268
rect 1942 252 1945 268
rect 1998 262 2001 298
rect 2006 252 2009 318
rect 2024 303 2026 307
rect 2030 303 2033 307
rect 2037 303 2040 307
rect 1846 162 1849 228
rect 1862 192 1865 208
rect 1742 152 1745 158
rect 1762 148 1766 151
rect 1814 142 1817 148
rect 1766 132 1769 138
rect 1766 112 1769 128
rect 1814 112 1817 138
rect 1766 92 1769 98
rect 1682 78 1686 81
rect 1686 62 1689 78
rect 1694 72 1697 78
rect 1702 42 1705 78
rect 1742 62 1745 78
rect 1774 42 1777 78
rect 1782 72 1785 108
rect 1814 92 1817 98
rect 1782 52 1785 68
rect 1822 62 1825 138
rect 1830 112 1833 148
rect 1862 142 1865 148
rect 1854 132 1857 138
rect 1334 -22 1345 -19
rect 1486 -18 1489 8
rect 1512 3 1514 7
rect 1518 3 1521 7
rect 1525 3 1528 7
rect 1542 -18 1545 8
rect 1598 -18 1601 8
rect 1782 -18 1785 48
rect 1798 41 1801 58
rect 1810 48 1814 51
rect 1822 41 1825 48
rect 1798 38 1825 41
rect 1830 42 1833 108
rect 1870 92 1873 198
rect 1878 162 1881 228
rect 1910 182 1913 238
rect 1958 232 1961 238
rect 1974 232 1977 238
rect 1982 232 1985 238
rect 1990 232 1993 238
rect 1942 192 1945 208
rect 1914 158 1918 161
rect 1942 152 1945 158
rect 2014 151 2017 278
rect 2054 262 2057 418
rect 2074 358 2078 361
rect 2062 262 2065 348
rect 2070 342 2073 348
rect 2094 342 2097 428
rect 2110 402 2113 478
rect 2118 412 2121 448
rect 2126 441 2129 548
rect 2134 542 2137 618
rect 2206 582 2209 678
rect 2222 662 2225 688
rect 2146 558 2150 561
rect 2158 552 2161 558
rect 2146 548 2150 551
rect 2166 542 2169 578
rect 2198 542 2201 547
rect 2214 542 2217 658
rect 2254 652 2257 659
rect 2262 492 2265 698
rect 2334 692 2337 708
rect 2366 702 2369 908
rect 2374 852 2377 868
rect 2382 862 2385 898
rect 2390 872 2393 888
rect 2414 852 2417 858
rect 2406 802 2409 818
rect 2422 792 2425 1018
rect 2434 988 2438 991
rect 2446 961 2449 1028
rect 2446 958 2454 961
rect 2446 942 2449 948
rect 2478 942 2481 1018
rect 2486 992 2489 1108
rect 2558 1102 2561 1128
rect 2526 1092 2529 1098
rect 2494 1062 2497 1088
rect 2546 1068 2550 1071
rect 2566 1061 2569 1218
rect 2574 1192 2577 1248
rect 2574 1172 2577 1188
rect 2582 1182 2585 1258
rect 2590 1252 2593 1258
rect 2598 1232 2601 1338
rect 2622 1332 2625 1338
rect 2646 1322 2649 1348
rect 2654 1332 2657 1338
rect 2606 1312 2609 1318
rect 2606 1262 2609 1298
rect 2670 1272 2673 1388
rect 2678 1342 2681 1358
rect 2686 1352 2689 1358
rect 2694 1352 2697 1598
rect 2702 1392 2705 1828
rect 2718 1782 2721 1818
rect 2766 1812 2769 1938
rect 2798 1932 2801 1948
rect 2814 1932 2817 1948
rect 2870 1942 2873 1948
rect 2850 1938 2854 1941
rect 2790 1922 2793 1928
rect 2778 1918 2782 1921
rect 2774 1852 2777 1868
rect 2790 1832 2793 1868
rect 2814 1832 2817 1878
rect 2822 1852 2825 1938
rect 2838 1892 2841 1928
rect 2854 1892 2857 1908
rect 2862 1882 2865 1918
rect 2870 1892 2873 1938
rect 2878 1932 2881 1938
rect 2910 1932 2913 1988
rect 2966 1982 2969 2028
rect 2990 1992 2993 1998
rect 2950 1962 2953 1968
rect 2918 1952 2921 1958
rect 2958 1952 2961 1958
rect 2922 1948 2926 1951
rect 2910 1912 2913 1928
rect 2918 1892 2921 1938
rect 2926 1892 2929 1938
rect 2942 1932 2945 1938
rect 2966 1912 2969 1948
rect 2974 1942 2977 1988
rect 3006 1952 3009 1958
rect 3014 1952 3017 1968
rect 2982 1932 2985 1938
rect 2990 1902 2993 1948
rect 3030 1932 3033 1968
rect 3054 1952 3057 2008
rect 3042 1938 3046 1941
rect 3014 1892 3017 1908
rect 3040 1903 3042 1907
rect 3046 1903 3049 1907
rect 3053 1903 3056 1907
rect 3062 1902 3065 2068
rect 3070 1972 3073 2058
rect 3078 2052 3081 2068
rect 3094 2062 3097 2068
rect 3110 2052 3113 2088
rect 3134 2062 3137 2068
rect 3142 2052 3145 2118
rect 3166 2092 3169 2128
rect 3182 2092 3185 2118
rect 3150 2072 3153 2078
rect 3198 2072 3201 2078
rect 3206 2061 3209 2118
rect 3214 2092 3217 2098
rect 3222 2081 3225 2148
rect 3230 2142 3233 2148
rect 3222 2078 3230 2081
rect 3198 2058 3209 2061
rect 3078 1941 3081 2048
rect 3182 2042 3185 2048
rect 3126 2032 3129 2038
rect 3086 1952 3089 2008
rect 3102 1942 3105 1948
rect 3078 1938 3089 1941
rect 3070 1932 3073 1938
rect 2890 1888 2894 1891
rect 3022 1882 3025 1898
rect 3086 1892 3089 1938
rect 3094 1882 3097 1938
rect 3110 1932 3113 1998
rect 3118 1992 3121 2018
rect 3126 1962 3129 1968
rect 3134 1952 3137 1988
rect 3142 1962 3145 2018
rect 3198 2002 3201 2058
rect 3222 2052 3225 2068
rect 3206 2042 3209 2048
rect 3142 1952 3145 1958
rect 3150 1942 3153 1978
rect 3162 1958 3166 1961
rect 3174 1942 3177 1978
rect 3194 1958 3198 1961
rect 3206 1952 3209 2038
rect 3238 2031 3241 2118
rect 3246 2082 3249 2148
rect 3310 2142 3313 2168
rect 3326 2162 3329 2178
rect 3338 2148 3342 2151
rect 3254 2091 3257 2138
rect 3262 2122 3265 2138
rect 3254 2088 3262 2091
rect 3262 2082 3265 2088
rect 3270 2072 3273 2138
rect 3350 2132 3353 2138
rect 3290 2128 3294 2131
rect 3302 2112 3305 2118
rect 3326 2072 3329 2108
rect 3358 2102 3361 2148
rect 3374 2132 3377 2148
rect 3382 2122 3385 2138
rect 3366 2082 3369 2118
rect 3390 2102 3393 2148
rect 3406 2132 3409 2158
rect 3414 2152 3417 2298
rect 3486 2282 3489 2548
rect 3510 2518 3518 2521
rect 3510 2482 3513 2518
rect 3510 2462 3513 2468
rect 3522 2458 3526 2461
rect 3494 2352 3497 2458
rect 3518 2392 3521 2448
rect 3534 2442 3537 2448
rect 3526 2361 3529 2418
rect 3518 2358 3529 2361
rect 3506 2348 3510 2351
rect 3430 2252 3433 2268
rect 3454 2262 3457 2268
rect 3494 2262 3497 2318
rect 3510 2252 3513 2258
rect 3450 2248 3454 2251
rect 3422 2222 3425 2228
rect 3422 2142 3425 2208
rect 3430 2202 3433 2248
rect 3470 2192 3473 2238
rect 3430 2152 3433 2158
rect 3438 2142 3441 2188
rect 3478 2142 3481 2198
rect 3458 2128 3462 2131
rect 3322 2068 3326 2071
rect 3378 2068 3382 2071
rect 3350 2062 3353 2068
rect 3322 2058 3326 2061
rect 3362 2058 3366 2061
rect 3354 2048 3358 2051
rect 3290 2038 3294 2041
rect 3230 2028 3241 2031
rect 3230 1992 3233 2028
rect 3238 2012 3241 2018
rect 3186 1948 3190 1951
rect 3230 1951 3233 1988
rect 3246 1962 3249 1968
rect 3266 1958 3270 1961
rect 3230 1948 3238 1951
rect 3266 1948 3270 1951
rect 3282 1948 3286 1951
rect 3294 1942 3297 1968
rect 3302 1952 3305 1958
rect 3358 1951 3361 1958
rect 3210 1938 3214 1941
rect 3306 1938 3310 1941
rect 3230 1932 3233 1938
rect 3238 1932 3241 1938
rect 3162 1928 3166 1931
rect 3118 1912 3121 1928
rect 3110 1908 3118 1911
rect 3110 1882 3113 1908
rect 3118 1882 3121 1888
rect 2846 1872 2849 1878
rect 2866 1868 2870 1871
rect 2830 1862 2833 1868
rect 2842 1858 2846 1861
rect 2758 1792 2761 1798
rect 2790 1792 2793 1798
rect 2798 1792 2801 1818
rect 2722 1768 2726 1771
rect 2718 1752 2721 1758
rect 2790 1752 2793 1768
rect 2810 1748 2814 1751
rect 2730 1738 2734 1741
rect 2750 1732 2753 1748
rect 2830 1732 2833 1758
rect 2838 1732 2841 1738
rect 2854 1732 2857 1828
rect 2878 1802 2881 1878
rect 2930 1868 2934 1871
rect 2994 1868 2998 1871
rect 3082 1868 3086 1871
rect 2902 1862 2905 1868
rect 2918 1852 2921 1868
rect 2942 1862 2945 1868
rect 3006 1862 3009 1868
rect 3074 1858 3078 1861
rect 2878 1752 2881 1798
rect 2894 1752 2897 1758
rect 2902 1752 2905 1818
rect 2918 1772 2921 1848
rect 2958 1842 2961 1848
rect 2934 1752 2937 1808
rect 2990 1792 2993 1858
rect 2998 1852 3001 1858
rect 3034 1848 3038 1851
rect 2882 1738 2886 1741
rect 2810 1728 2814 1731
rect 2710 1692 2713 1708
rect 2742 1702 2745 1718
rect 2774 1712 2777 1718
rect 2782 1702 2785 1728
rect 2718 1672 2721 1678
rect 2726 1662 2729 1668
rect 2750 1662 2753 1668
rect 2782 1662 2785 1668
rect 2770 1658 2774 1661
rect 2738 1648 2742 1651
rect 2710 1542 2713 1548
rect 2718 1512 2721 1548
rect 2726 1502 2729 1618
rect 2750 1592 2753 1608
rect 2774 1592 2777 1628
rect 2798 1602 2801 1718
rect 2822 1682 2825 1718
rect 2810 1658 2814 1661
rect 2842 1658 2846 1661
rect 2738 1568 2742 1571
rect 2738 1558 2742 1561
rect 2750 1552 2753 1558
rect 2790 1532 2793 1538
rect 2798 1532 2801 1588
rect 2806 1572 2809 1578
rect 2822 1551 2825 1618
rect 2814 1548 2825 1551
rect 2830 1562 2833 1638
rect 2878 1632 2881 1658
rect 2894 1642 2897 1648
rect 2854 1582 2857 1588
rect 2838 1562 2841 1568
rect 2830 1552 2833 1558
rect 2862 1552 2865 1618
rect 2902 1592 2905 1748
rect 2910 1692 2913 1718
rect 2910 1652 2913 1668
rect 2918 1632 2921 1718
rect 2934 1672 2937 1748
rect 2942 1742 2945 1778
rect 2962 1748 2966 1751
rect 2998 1742 3001 1838
rect 3094 1812 3097 1878
rect 3142 1872 3145 1888
rect 3222 1882 3225 1918
rect 3230 1882 3233 1898
rect 3270 1872 3273 1938
rect 3314 1928 3318 1931
rect 3326 1892 3329 1948
rect 3106 1858 3110 1861
rect 3118 1852 3121 1858
rect 3090 1758 3094 1761
rect 3030 1752 3033 1758
rect 3066 1748 3070 1751
rect 3066 1738 3070 1741
rect 2942 1732 2945 1738
rect 2950 1672 2953 1718
rect 2966 1711 2969 1728
rect 2974 1722 2977 1738
rect 3086 1732 3089 1738
rect 2966 1708 2977 1711
rect 2966 1682 2969 1688
rect 2926 1652 2929 1658
rect 2870 1552 2873 1568
rect 2878 1562 2881 1568
rect 2894 1562 2897 1568
rect 2850 1548 2854 1551
rect 2734 1522 2737 1528
rect 2806 1522 2809 1528
rect 2726 1482 2729 1488
rect 2758 1482 2761 1508
rect 2798 1472 2801 1478
rect 2738 1468 2742 1471
rect 2710 1462 2713 1468
rect 2762 1458 2766 1461
rect 2778 1458 2782 1461
rect 2722 1448 2726 1451
rect 2770 1448 2774 1451
rect 2814 1422 2817 1548
rect 2822 1532 2825 1538
rect 2862 1532 2865 1538
rect 2878 1492 2881 1548
rect 2926 1542 2929 1648
rect 2934 1542 2937 1658
rect 2942 1652 2945 1668
rect 2958 1652 2961 1658
rect 2950 1552 2953 1558
rect 2958 1552 2961 1648
rect 2974 1582 2977 1708
rect 2998 1681 3001 1728
rect 3078 1712 3081 1718
rect 3040 1703 3042 1707
rect 3046 1703 3049 1707
rect 3053 1703 3056 1707
rect 3094 1702 3097 1718
rect 3010 1688 3014 1691
rect 3062 1682 3065 1688
rect 3102 1682 3105 1818
rect 3142 1811 3145 1858
rect 3150 1822 3153 1868
rect 3162 1848 3166 1851
rect 3174 1842 3177 1868
rect 3222 1862 3225 1868
rect 3234 1858 3238 1861
rect 3206 1852 3209 1858
rect 3246 1822 3249 1868
rect 3254 1852 3257 1858
rect 3262 1852 3265 1858
rect 3278 1822 3281 1858
rect 3286 1852 3289 1868
rect 3318 1863 3321 1878
rect 3342 1862 3345 1938
rect 3382 1932 3385 2068
rect 3398 2022 3401 2078
rect 3430 2052 3433 2059
rect 3430 1962 3433 1968
rect 3418 1958 3422 1961
rect 3390 1952 3393 1958
rect 3446 1952 3449 2068
rect 3462 2062 3465 2068
rect 3470 1992 3473 2008
rect 3486 1992 3489 2138
rect 3518 2082 3521 2358
rect 3526 2332 3529 2348
rect 3558 2342 3561 2348
rect 3526 2302 3529 2328
rect 3550 2292 3553 2298
rect 3558 2272 3561 2298
rect 3542 2192 3545 2248
rect 3542 2062 3545 2118
rect 3466 1968 3470 1971
rect 3482 1968 3486 1971
rect 3386 1928 3393 1931
rect 3378 1888 3382 1891
rect 3390 1872 3393 1928
rect 3446 1882 3449 1948
rect 3454 1942 3457 1948
rect 3478 1942 3481 1948
rect 3454 1872 3457 1938
rect 3478 1892 3481 1938
rect 3494 1932 3497 2018
rect 3502 2012 3505 2058
rect 3526 2022 3529 2058
rect 3558 2042 3561 2048
rect 3502 1952 3505 1958
rect 3510 1902 3513 2018
rect 3518 1972 3521 1978
rect 3522 1948 3526 1951
rect 3558 1942 3561 1948
rect 3518 1892 3521 1938
rect 3510 1882 3513 1888
rect 3142 1808 3153 1811
rect 3150 1792 3153 1808
rect 3158 1761 3161 1818
rect 3278 1792 3281 1818
rect 3230 1782 3233 1788
rect 3286 1782 3289 1848
rect 3294 1762 3297 1788
rect 3366 1782 3369 1788
rect 3358 1762 3361 1778
rect 3158 1758 3166 1761
rect 3258 1758 3262 1761
rect 3390 1761 3393 1868
rect 3398 1862 3401 1868
rect 3410 1858 3414 1861
rect 3450 1859 3454 1862
rect 3526 1862 3529 1878
rect 3410 1848 3414 1851
rect 3398 1792 3401 1848
rect 3558 1842 3561 1848
rect 3386 1758 3393 1761
rect 3110 1752 3113 1758
rect 3130 1728 3134 1731
rect 3110 1682 3113 1728
rect 3142 1712 3145 1738
rect 3150 1732 3153 1748
rect 3182 1742 3185 1758
rect 3206 1752 3209 1758
rect 3258 1748 3262 1751
rect 3302 1742 3305 1758
rect 3354 1748 3358 1751
rect 3374 1742 3377 1748
rect 3226 1738 3230 1741
rect 3266 1738 3270 1741
rect 3298 1738 3302 1741
rect 3206 1732 3209 1738
rect 3238 1732 3241 1738
rect 3162 1688 3166 1691
rect 3174 1682 3177 1688
rect 2998 1678 3006 1681
rect 3034 1678 3038 1681
rect 2982 1672 2985 1678
rect 3102 1662 3105 1678
rect 3150 1662 3153 1678
rect 3074 1658 3078 1661
rect 3146 1658 3150 1661
rect 2990 1592 2993 1598
rect 2998 1592 3001 1618
rect 2994 1568 2998 1571
rect 2910 1532 2913 1538
rect 2942 1531 2945 1538
rect 2938 1528 2945 1531
rect 2886 1492 2889 1528
rect 2918 1512 2921 1528
rect 2926 1522 2929 1528
rect 2822 1482 2825 1488
rect 2902 1482 2905 1488
rect 2866 1478 2870 1481
rect 2878 1478 2886 1481
rect 2846 1472 2849 1478
rect 2866 1468 2870 1471
rect 2834 1458 2838 1461
rect 2850 1458 2854 1461
rect 2782 1372 2785 1418
rect 2838 1392 2841 1448
rect 2862 1402 2865 1418
rect 2862 1392 2865 1398
rect 2726 1362 2729 1368
rect 2842 1358 2846 1361
rect 2702 1352 2705 1358
rect 2766 1352 2769 1358
rect 2754 1348 2758 1351
rect 2710 1332 2713 1338
rect 2682 1328 2686 1331
rect 2618 1268 2622 1271
rect 2650 1268 2654 1271
rect 2698 1268 2702 1271
rect 2618 1248 2622 1251
rect 2582 1152 2585 1168
rect 2606 1142 2609 1228
rect 2630 1212 2633 1258
rect 2638 1242 2641 1248
rect 2614 1152 2617 1168
rect 2562 1058 2569 1061
rect 2536 1003 2538 1007
rect 2542 1003 2545 1007
rect 2549 1003 2552 1007
rect 2558 972 2561 1018
rect 2574 952 2577 1138
rect 2618 1078 2622 1081
rect 2630 1072 2633 1198
rect 2646 1181 2649 1218
rect 2642 1178 2649 1181
rect 2654 1171 2657 1248
rect 2646 1168 2657 1171
rect 2646 1152 2649 1168
rect 2662 1142 2665 1218
rect 2678 1152 2681 1158
rect 2694 1142 2697 1268
rect 2710 1192 2713 1328
rect 2718 1322 2721 1348
rect 2726 1342 2729 1348
rect 2738 1338 2742 1341
rect 2754 1338 2758 1341
rect 2782 1312 2785 1358
rect 2790 1292 2793 1358
rect 2878 1352 2881 1478
rect 2886 1462 2889 1468
rect 2902 1462 2905 1478
rect 2910 1462 2913 1468
rect 2918 1462 2921 1508
rect 2926 1462 2929 1468
rect 2934 1432 2937 1508
rect 2942 1492 2945 1518
rect 2950 1512 2953 1538
rect 2974 1522 2977 1528
rect 2942 1482 2945 1488
rect 2950 1462 2953 1498
rect 2966 1482 2969 1518
rect 2974 1472 2977 1478
rect 2982 1472 2985 1558
rect 3030 1552 3033 1658
rect 3086 1652 3089 1658
rect 3134 1652 3137 1658
rect 3190 1652 3193 1718
rect 3198 1712 3201 1728
rect 3214 1682 3217 1688
rect 3050 1648 3054 1651
rect 3178 1648 3182 1651
rect 3198 1642 3201 1668
rect 3246 1662 3249 1678
rect 3262 1672 3265 1678
rect 3274 1668 3278 1671
rect 3254 1662 3257 1668
rect 3210 1658 3214 1661
rect 3122 1618 3126 1621
rect 3070 1552 3073 1618
rect 3086 1612 3089 1618
rect 3134 1612 3137 1618
rect 3078 1552 3081 1558
rect 3010 1548 3014 1551
rect 2990 1542 2993 1548
rect 3070 1532 3073 1538
rect 3030 1522 3033 1528
rect 2958 1452 2961 1468
rect 2990 1462 2993 1488
rect 2998 1471 3001 1518
rect 3022 1502 3025 1518
rect 3040 1503 3042 1507
rect 3046 1503 3049 1507
rect 3053 1503 3056 1507
rect 3010 1478 3014 1481
rect 3022 1472 3025 1478
rect 3054 1472 3057 1478
rect 2998 1468 3006 1471
rect 3034 1468 3038 1471
rect 2970 1458 2974 1461
rect 3030 1452 3033 1458
rect 2990 1432 2993 1448
rect 3062 1442 3065 1448
rect 2910 1392 2913 1408
rect 2890 1378 2894 1381
rect 2926 1362 2929 1418
rect 2826 1348 2830 1351
rect 2866 1348 2870 1351
rect 2814 1342 2817 1348
rect 2926 1342 2929 1348
rect 2934 1342 2937 1428
rect 2994 1378 2998 1381
rect 2978 1358 2982 1361
rect 2942 1342 2945 1358
rect 2954 1348 2958 1351
rect 2966 1342 2969 1358
rect 2986 1348 2990 1351
rect 2998 1342 3001 1348
rect 3006 1342 3009 1348
rect 2802 1338 2806 1341
rect 2822 1332 2825 1338
rect 2958 1332 2961 1338
rect 2842 1328 2846 1331
rect 2854 1322 2857 1328
rect 2758 1272 2761 1278
rect 2782 1262 2785 1268
rect 2738 1258 2742 1261
rect 2718 1252 2721 1258
rect 2770 1248 2774 1251
rect 2702 1142 2705 1148
rect 2710 1142 2713 1148
rect 2718 1142 2721 1168
rect 2726 1152 2729 1248
rect 2746 1238 2750 1241
rect 2798 1222 2801 1318
rect 2830 1282 2833 1298
rect 2846 1292 2849 1298
rect 2942 1292 2945 1318
rect 2990 1292 2993 1318
rect 3014 1292 3017 1298
rect 2878 1278 2894 1281
rect 2814 1232 2817 1258
rect 2834 1248 2838 1251
rect 2742 1142 2745 1158
rect 2750 1142 2753 1218
rect 2782 1152 2785 1178
rect 2766 1141 2769 1148
rect 2790 1142 2793 1168
rect 2846 1162 2849 1268
rect 2854 1262 2857 1268
rect 2878 1252 2881 1278
rect 2918 1272 2921 1278
rect 2966 1272 2969 1278
rect 2998 1272 3001 1278
rect 2890 1268 2894 1271
rect 3010 1268 3014 1271
rect 2974 1262 2977 1268
rect 2898 1258 2902 1261
rect 2914 1258 2918 1261
rect 2886 1252 2889 1258
rect 2802 1148 2806 1151
rect 2766 1138 2785 1141
rect 2814 1141 2817 1158
rect 2862 1152 2865 1248
rect 2926 1242 2929 1258
rect 2942 1252 2945 1258
rect 3014 1252 3017 1258
rect 2954 1248 2958 1251
rect 2918 1192 2921 1218
rect 2942 1192 2945 1198
rect 2966 1192 2969 1238
rect 3022 1212 3025 1438
rect 3054 1422 3057 1428
rect 3062 1392 3065 1438
rect 3030 1352 3033 1368
rect 3070 1332 3073 1468
rect 3086 1362 3089 1608
rect 3150 1592 3153 1638
rect 3190 1622 3193 1628
rect 3190 1592 3193 1608
rect 3154 1568 3158 1571
rect 3118 1552 3121 1568
rect 3142 1562 3145 1568
rect 3174 1562 3177 1568
rect 3166 1552 3169 1558
rect 3126 1542 3129 1548
rect 3182 1542 3185 1588
rect 3206 1552 3209 1638
rect 3230 1612 3233 1618
rect 3230 1552 3233 1608
rect 3278 1562 3281 1618
rect 3286 1552 3289 1728
rect 3302 1672 3305 1718
rect 3326 1682 3329 1688
rect 3314 1678 3318 1681
rect 3342 1672 3345 1678
rect 3294 1662 3297 1668
rect 3342 1652 3345 1658
rect 3322 1648 3326 1651
rect 3350 1592 3353 1738
rect 3382 1692 3385 1758
rect 3358 1672 3361 1678
rect 3370 1668 3374 1671
rect 3358 1642 3361 1668
rect 3366 1652 3369 1658
rect 3374 1592 3377 1658
rect 3382 1642 3385 1668
rect 3398 1662 3401 1748
rect 3406 1742 3409 1778
rect 3418 1738 3422 1741
rect 3414 1672 3417 1698
rect 3438 1692 3441 1818
rect 3470 1722 3473 1728
rect 3454 1682 3457 1688
rect 3430 1672 3433 1678
rect 3426 1658 3430 1661
rect 3394 1648 3398 1651
rect 3414 1651 3417 1658
rect 3414 1648 3425 1651
rect 3406 1642 3409 1648
rect 3334 1562 3337 1568
rect 3422 1562 3425 1648
rect 3394 1558 3398 1561
rect 3366 1552 3369 1558
rect 3354 1548 3358 1551
rect 3410 1548 3414 1551
rect 3102 1522 3105 1528
rect 3106 1459 3110 1462
rect 3134 1462 3137 1538
rect 3146 1528 3150 1531
rect 3206 1512 3209 1548
rect 3226 1538 3230 1541
rect 3214 1532 3217 1538
rect 3230 1522 3233 1528
rect 3166 1482 3169 1488
rect 3222 1471 3225 1518
rect 3270 1512 3273 1548
rect 3370 1538 3414 1541
rect 3330 1518 3334 1521
rect 3302 1492 3305 1508
rect 3274 1478 3278 1481
rect 3290 1478 3305 1481
rect 3222 1468 3230 1471
rect 3254 1468 3281 1471
rect 3238 1462 3241 1468
rect 3254 1462 3257 1468
rect 3178 1458 3182 1461
rect 3266 1458 3270 1461
rect 3278 1461 3281 1468
rect 3302 1471 3305 1478
rect 3302 1468 3326 1471
rect 3294 1462 3297 1468
rect 3278 1458 3286 1461
rect 3322 1458 3329 1461
rect 3170 1448 3174 1451
rect 3190 1442 3193 1458
rect 3222 1452 3225 1458
rect 3230 1452 3233 1458
rect 3198 1448 3206 1451
rect 3102 1392 3105 1398
rect 3150 1392 3153 1438
rect 3078 1342 3081 1348
rect 3086 1342 3089 1348
rect 3166 1342 3169 1348
rect 3114 1338 3118 1341
rect 3174 1332 3177 1338
rect 3040 1303 3042 1307
rect 3046 1303 3049 1307
rect 3053 1303 3056 1307
rect 3086 1292 3089 1298
rect 3150 1272 3153 1278
rect 3034 1268 3038 1271
rect 3106 1268 3110 1271
rect 3054 1262 3057 1268
rect 3114 1258 3118 1261
rect 3126 1232 3129 1248
rect 3150 1242 3153 1268
rect 3014 1192 3017 1198
rect 3070 1192 3073 1208
rect 3158 1192 3161 1268
rect 3166 1262 3169 1268
rect 3174 1251 3177 1328
rect 3190 1312 3193 1338
rect 3198 1322 3201 1448
rect 3246 1432 3249 1458
rect 3326 1452 3329 1458
rect 3270 1442 3273 1448
rect 3318 1392 3321 1438
rect 3342 1422 3345 1538
rect 3422 1522 3425 1558
rect 3438 1552 3441 1678
rect 3446 1652 3449 1678
rect 3478 1672 3481 1788
rect 3494 1752 3497 1798
rect 3486 1712 3489 1738
rect 3502 1711 3505 1808
rect 3510 1762 3513 1828
rect 3538 1748 3542 1751
rect 3530 1738 3534 1741
rect 3558 1732 3561 1738
rect 3514 1728 3518 1731
rect 3514 1718 3518 1721
rect 3502 1708 3513 1711
rect 3454 1662 3457 1668
rect 3470 1662 3473 1668
rect 3478 1572 3481 1668
rect 3486 1662 3489 1698
rect 3510 1692 3513 1708
rect 3526 1702 3529 1718
rect 3502 1682 3505 1688
rect 3530 1678 3534 1681
rect 3486 1632 3489 1658
rect 3498 1648 3502 1651
rect 3478 1552 3481 1558
rect 3430 1548 3438 1551
rect 3350 1472 3353 1518
rect 3382 1492 3385 1508
rect 3398 1492 3401 1498
rect 3362 1478 3374 1481
rect 3394 1478 3398 1481
rect 3430 1472 3433 1548
rect 3442 1538 3446 1541
rect 3466 1538 3470 1541
rect 3454 1501 3457 1528
rect 3462 1511 3465 1518
rect 3462 1508 3470 1511
rect 3454 1498 3465 1501
rect 3402 1468 3406 1471
rect 3350 1442 3353 1468
rect 3366 1432 3369 1468
rect 3414 1462 3417 1468
rect 3438 1462 3441 1478
rect 3446 1472 3449 1498
rect 3454 1472 3457 1478
rect 3418 1448 3422 1451
rect 3382 1431 3385 1448
rect 3374 1428 3385 1431
rect 3206 1362 3209 1388
rect 3274 1368 3278 1371
rect 3286 1352 3289 1358
rect 3226 1348 3230 1351
rect 3242 1348 3249 1351
rect 3234 1338 3238 1341
rect 3194 1278 3198 1281
rect 3206 1272 3209 1318
rect 3214 1292 3217 1318
rect 3238 1272 3241 1338
rect 3246 1332 3249 1348
rect 3278 1342 3281 1348
rect 3334 1342 3337 1388
rect 3342 1352 3345 1398
rect 3314 1328 3318 1331
rect 3254 1302 3257 1328
rect 3254 1282 3257 1288
rect 3270 1262 3273 1288
rect 3278 1262 3281 1268
rect 3166 1248 3177 1251
rect 3182 1252 3185 1258
rect 3190 1252 3193 1258
rect 3202 1248 3206 1251
rect 2870 1182 2873 1188
rect 3026 1158 3030 1161
rect 2798 1138 2817 1141
rect 2638 1072 2641 1138
rect 2662 1122 2665 1128
rect 2654 1072 2657 1078
rect 2678 1072 2681 1138
rect 2694 1092 2697 1118
rect 2702 1082 2705 1138
rect 2762 1128 2766 1131
rect 2782 1131 2785 1138
rect 2798 1131 2801 1138
rect 2782 1128 2801 1131
rect 2822 1132 2825 1138
rect 2718 1092 2721 1128
rect 2734 1102 2737 1128
rect 2774 1078 2777 1128
rect 2686 1072 2689 1078
rect 2610 1068 2614 1071
rect 2602 1058 2609 1061
rect 2606 1052 2609 1058
rect 2590 992 2593 1038
rect 2538 948 2542 951
rect 2602 948 2606 951
rect 2466 938 2470 941
rect 2430 872 2433 888
rect 2438 862 2441 938
rect 2462 892 2465 918
rect 2454 882 2457 888
rect 2466 878 2470 881
rect 2446 872 2449 878
rect 2502 872 2505 918
rect 2510 872 2513 918
rect 2522 878 2526 881
rect 2498 858 2502 861
rect 2486 852 2489 858
rect 2518 852 2521 858
rect 2498 848 2502 851
rect 2474 838 2478 841
rect 2550 822 2553 918
rect 2614 872 2617 978
rect 2622 892 2625 918
rect 2602 868 2606 871
rect 2578 858 2582 861
rect 2590 832 2593 838
rect 2486 792 2489 818
rect 2536 803 2538 807
rect 2542 803 2545 807
rect 2549 803 2552 807
rect 2406 752 2409 788
rect 2426 758 2430 761
rect 2450 758 2454 761
rect 2414 752 2417 758
rect 2498 748 2502 751
rect 2534 751 2537 758
rect 2374 712 2377 748
rect 2438 742 2441 748
rect 2462 742 2465 748
rect 2470 742 2473 748
rect 2550 742 2553 748
rect 2454 732 2457 738
rect 2426 728 2430 731
rect 2490 728 2494 731
rect 2402 718 2406 721
rect 2542 712 2545 738
rect 2558 712 2561 818
rect 2606 771 2609 788
rect 2602 768 2609 771
rect 2606 752 2609 768
rect 2322 688 2326 691
rect 2350 682 2353 688
rect 2338 678 2342 681
rect 2370 668 2374 671
rect 2286 662 2289 668
rect 2326 652 2329 658
rect 2366 652 2369 658
rect 2286 572 2289 638
rect 2274 558 2278 561
rect 2286 552 2289 568
rect 2310 552 2313 558
rect 2318 552 2321 578
rect 2326 552 2329 648
rect 2382 642 2385 658
rect 2390 652 2393 658
rect 2398 652 2401 678
rect 2414 672 2417 678
rect 2406 662 2409 668
rect 2366 572 2369 618
rect 2374 592 2377 608
rect 2346 558 2350 561
rect 2362 548 2366 551
rect 2358 542 2361 548
rect 2298 538 2302 541
rect 2310 532 2313 538
rect 2270 502 2273 528
rect 2294 488 2310 491
rect 2142 472 2145 488
rect 2174 472 2177 478
rect 2186 468 2190 471
rect 2134 452 2137 468
rect 2230 462 2233 468
rect 2126 438 2137 441
rect 2134 392 2137 438
rect 2142 422 2145 458
rect 2150 442 2153 448
rect 2166 442 2169 448
rect 2174 432 2177 458
rect 2102 352 2105 378
rect 2134 368 2142 371
rect 2106 338 2110 341
rect 2078 332 2081 338
rect 2122 328 2126 331
rect 2134 321 2137 368
rect 2146 348 2150 351
rect 2126 318 2137 321
rect 2090 278 2094 281
rect 2098 268 2102 271
rect 2026 258 2030 261
rect 2066 258 2070 261
rect 2022 162 2025 258
rect 2050 248 2054 251
rect 2066 248 2070 251
rect 2034 228 2038 231
rect 2054 171 2057 248
rect 2078 222 2081 268
rect 2110 262 2113 268
rect 2118 261 2121 318
rect 2126 272 2129 318
rect 2158 312 2161 358
rect 2166 332 2169 428
rect 2182 362 2185 458
rect 2238 452 2241 478
rect 2254 472 2257 478
rect 2250 468 2254 471
rect 2294 462 2297 488
rect 2342 481 2345 518
rect 2374 492 2377 578
rect 2386 548 2390 551
rect 2390 512 2393 528
rect 2406 492 2409 638
rect 2430 582 2433 678
rect 2438 672 2441 678
rect 2494 672 2497 688
rect 2438 658 2446 661
rect 2474 658 2478 661
rect 2438 652 2441 658
rect 2466 648 2470 651
rect 2510 642 2513 678
rect 2542 672 2545 708
rect 2466 638 2470 641
rect 2542 622 2545 668
rect 2558 652 2561 659
rect 2446 552 2449 558
rect 2430 492 2433 528
rect 2342 478 2350 481
rect 2302 472 2305 478
rect 2318 462 2321 478
rect 2334 472 2337 478
rect 2398 472 2401 478
rect 2454 472 2457 548
rect 2478 542 2481 618
rect 2536 603 2538 607
rect 2542 603 2545 607
rect 2549 603 2552 607
rect 2558 582 2561 598
rect 2566 592 2569 748
rect 2614 742 2617 818
rect 2630 772 2633 1068
rect 2662 1062 2665 1068
rect 2682 1058 2686 1061
rect 2638 992 2641 1058
rect 2638 952 2641 988
rect 2646 822 2649 1058
rect 2702 1012 2705 1068
rect 2710 1052 2713 1058
rect 2718 1052 2721 1078
rect 2798 1072 2801 1108
rect 2806 1092 2809 1098
rect 2734 1052 2737 1058
rect 2742 1042 2745 1068
rect 2718 992 2721 1008
rect 2750 982 2753 1068
rect 2766 1042 2769 1058
rect 2782 1042 2785 1058
rect 2798 1042 2801 1068
rect 2806 1062 2809 1068
rect 2806 1032 2809 1048
rect 2814 1032 2817 1118
rect 2830 1112 2833 1148
rect 2834 1078 2838 1081
rect 2846 1072 2849 1078
rect 2846 1052 2849 1058
rect 2862 1051 2865 1148
rect 2882 1138 2886 1141
rect 2902 1132 2905 1158
rect 2878 1072 2881 1118
rect 2894 1112 2897 1128
rect 2902 1092 2905 1098
rect 2910 1072 2913 1078
rect 2890 1068 2894 1071
rect 2878 1062 2881 1068
rect 2858 1048 2865 1051
rect 2918 1061 2921 1148
rect 2926 1082 2929 1138
rect 2934 1072 2937 1138
rect 2950 1132 2953 1148
rect 2962 1138 2966 1141
rect 2982 1092 2985 1158
rect 2994 1138 2998 1141
rect 2994 1128 2998 1131
rect 2930 1068 2934 1071
rect 2910 1058 2921 1061
rect 2938 1058 2942 1061
rect 2954 1058 2958 1061
rect 2870 1052 2873 1058
rect 2774 952 2777 958
rect 2806 952 2809 958
rect 2722 948 2726 951
rect 2662 942 2665 948
rect 2654 852 2657 938
rect 2710 932 2713 938
rect 2734 932 2737 948
rect 2742 932 2745 938
rect 2694 902 2697 918
rect 2774 912 2777 938
rect 2710 892 2713 908
rect 2742 892 2745 908
rect 2738 878 2742 881
rect 2750 872 2753 878
rect 2674 868 2678 871
rect 2674 858 2678 861
rect 2678 812 2681 848
rect 2694 842 2697 848
rect 2710 822 2713 848
rect 2750 822 2753 858
rect 2678 792 2681 808
rect 2642 778 2646 781
rect 2626 748 2630 751
rect 2606 732 2609 738
rect 2614 722 2617 738
rect 2622 732 2625 738
rect 2630 732 2633 738
rect 2638 692 2641 758
rect 2654 742 2657 758
rect 2742 752 2745 768
rect 2710 742 2713 748
rect 2662 732 2665 738
rect 2722 728 2726 731
rect 2654 682 2657 688
rect 2662 682 2665 688
rect 2710 682 2713 688
rect 2726 682 2729 718
rect 2734 712 2737 748
rect 2746 738 2750 741
rect 2742 682 2745 718
rect 2758 692 2761 888
rect 2766 872 2769 878
rect 2766 752 2769 868
rect 2774 842 2777 868
rect 2782 862 2785 948
rect 2798 922 2801 928
rect 2798 882 2801 918
rect 2806 892 2809 948
rect 2822 892 2825 1008
rect 2830 992 2833 998
rect 2846 992 2849 1008
rect 2858 958 2862 961
rect 2866 958 2873 961
rect 2830 932 2833 938
rect 2846 932 2849 948
rect 2870 932 2873 958
rect 2814 882 2817 888
rect 2830 882 2833 928
rect 2846 892 2849 928
rect 2878 912 2881 1058
rect 2902 972 2905 1048
rect 2894 942 2897 948
rect 2910 942 2913 1058
rect 2938 1048 2942 1051
rect 2918 982 2921 1018
rect 2942 1012 2945 1028
rect 2950 1012 2953 1048
rect 2974 1012 2977 1078
rect 2998 1072 3001 1108
rect 3006 1102 3009 1138
rect 3014 1132 3017 1148
rect 3030 1128 3038 1131
rect 3006 1082 3009 1098
rect 2990 1062 2993 1068
rect 2998 1062 3001 1068
rect 3014 1002 3017 1128
rect 3030 1102 3033 1128
rect 3040 1103 3042 1107
rect 3046 1103 3049 1107
rect 3053 1103 3056 1107
rect 3022 1032 3025 1058
rect 3046 1032 3049 1078
rect 3062 1072 3065 1188
rect 3086 1151 3089 1168
rect 3086 1148 3094 1151
rect 3106 1148 3110 1151
rect 3078 1132 3081 1148
rect 3062 1052 3065 1058
rect 2918 932 2921 958
rect 2934 952 2937 958
rect 2942 952 2945 978
rect 2962 958 2966 961
rect 2978 948 2982 951
rect 2926 941 2929 948
rect 2998 942 3001 948
rect 3046 942 3049 988
rect 3054 942 3057 948
rect 2926 938 2934 941
rect 2978 938 2982 941
rect 2950 922 2953 928
rect 2790 872 2793 878
rect 2854 872 2857 878
rect 2862 862 2865 908
rect 2958 902 2961 928
rect 2966 892 2969 928
rect 2902 862 2905 878
rect 2926 872 2929 878
rect 2942 872 2945 888
rect 2974 872 2977 898
rect 2966 868 2974 871
rect 2866 858 2870 861
rect 2806 822 2809 848
rect 2830 822 2833 858
rect 2838 852 2841 858
rect 2926 852 2929 858
rect 2882 848 2886 851
rect 2914 848 2918 851
rect 2782 802 2785 818
rect 2786 768 2790 771
rect 2798 752 2801 788
rect 2774 742 2777 748
rect 2794 738 2798 741
rect 2626 678 2630 681
rect 2694 672 2697 678
rect 2766 672 2769 728
rect 2646 662 2649 668
rect 2626 638 2630 641
rect 2670 622 2673 668
rect 2678 662 2681 668
rect 2686 652 2689 658
rect 2742 652 2745 659
rect 2706 648 2710 651
rect 2774 642 2777 728
rect 2806 722 2809 748
rect 2822 732 2825 758
rect 2838 741 2841 848
rect 2886 822 2889 848
rect 2934 842 2937 858
rect 2950 812 2953 868
rect 2966 852 2969 868
rect 2982 862 2985 908
rect 2990 892 2993 938
rect 3040 903 3042 907
rect 3046 903 3049 907
rect 3053 903 3056 907
rect 3030 862 3033 878
rect 3038 872 3041 888
rect 3022 851 3025 858
rect 3046 851 3049 858
rect 3022 848 3049 851
rect 2954 778 2958 781
rect 2846 752 2849 758
rect 2854 752 2857 778
rect 2890 747 2894 750
rect 2958 742 2961 748
rect 2838 738 2849 741
rect 2622 592 2625 608
rect 2654 572 2657 578
rect 2602 558 2606 561
rect 2582 552 2585 558
rect 2514 548 2518 551
rect 2614 548 2622 551
rect 2498 538 2502 541
rect 2546 538 2550 541
rect 2494 522 2497 528
rect 2486 492 2489 508
rect 2510 502 2513 538
rect 2518 528 2526 531
rect 2570 528 2574 531
rect 2426 468 2430 471
rect 2246 452 2249 458
rect 2302 452 2305 458
rect 2310 452 2313 458
rect 2206 382 2209 418
rect 2246 412 2249 448
rect 2230 392 2233 398
rect 2278 362 2281 448
rect 2302 392 2305 428
rect 2210 358 2214 361
rect 2250 358 2254 361
rect 2182 352 2185 358
rect 2318 352 2321 438
rect 2326 412 2329 458
rect 2334 452 2337 468
rect 2342 462 2345 468
rect 2350 462 2353 468
rect 2454 462 2457 468
rect 2378 458 2385 461
rect 2366 412 2369 448
rect 2374 442 2377 448
rect 2350 392 2353 408
rect 2358 362 2361 378
rect 2194 348 2198 351
rect 2242 348 2246 351
rect 2174 342 2177 348
rect 2206 342 2209 348
rect 2190 332 2193 338
rect 2166 302 2169 328
rect 2222 322 2225 338
rect 2266 328 2270 331
rect 2278 322 2281 348
rect 2306 338 2310 341
rect 2326 332 2329 338
rect 2306 328 2310 331
rect 2150 272 2153 298
rect 2254 292 2257 308
rect 2334 292 2337 358
rect 2366 352 2369 398
rect 2382 352 2385 458
rect 2390 422 2393 458
rect 2406 352 2409 448
rect 2430 442 2433 448
rect 2430 362 2433 438
rect 2446 422 2449 458
rect 2454 432 2457 458
rect 2494 451 2497 468
rect 2490 448 2497 451
rect 2502 452 2505 458
rect 2454 382 2457 388
rect 2346 328 2353 331
rect 2286 282 2289 288
rect 2290 278 2294 281
rect 2198 272 2201 278
rect 2326 272 2329 278
rect 2342 272 2345 298
rect 2210 268 2214 271
rect 2134 262 2137 268
rect 2222 262 2225 268
rect 2118 258 2129 261
rect 2146 258 2150 261
rect 2258 258 2262 261
rect 2054 168 2065 171
rect 2050 158 2054 161
rect 2062 152 2065 168
rect 2078 152 2081 158
rect 2010 148 2017 151
rect 2042 148 2046 151
rect 1886 132 1889 138
rect 1910 132 1913 138
rect 1926 122 1929 128
rect 1874 78 1878 81
rect 1902 81 1905 118
rect 1934 92 1937 128
rect 1942 112 1945 138
rect 1898 78 1905 81
rect 1910 78 1918 81
rect 1922 78 1926 81
rect 1846 72 1849 78
rect 1886 71 1889 78
rect 1886 68 1894 71
rect 1910 71 1913 78
rect 1902 68 1913 71
rect 1918 72 1921 78
rect 1942 72 1945 98
rect 1838 52 1841 68
rect 1902 61 1905 68
rect 1950 62 1953 148
rect 2006 142 2009 148
rect 2086 142 2089 258
rect 2094 252 2097 258
rect 2114 248 2118 251
rect 2126 232 2129 258
rect 2238 252 2241 258
rect 2270 252 2273 268
rect 2206 242 2209 248
rect 2254 242 2257 248
rect 2286 242 2289 248
rect 2130 158 2134 161
rect 2142 152 2145 158
rect 2158 152 2161 228
rect 2166 152 2169 178
rect 2222 152 2225 238
rect 2294 222 2297 268
rect 2302 262 2305 268
rect 2318 262 2321 268
rect 2318 232 2321 248
rect 2278 192 2281 198
rect 2258 158 2262 161
rect 2114 148 2118 151
rect 2210 148 2214 151
rect 2266 148 2278 151
rect 2118 142 2121 148
rect 2190 142 2193 148
rect 2286 142 2289 218
rect 2334 192 2337 228
rect 2342 182 2345 268
rect 2350 262 2353 328
rect 2374 312 2377 348
rect 2394 338 2398 341
rect 2382 331 2385 338
rect 2414 332 2417 358
rect 2422 342 2425 348
rect 2430 342 2433 348
rect 2382 328 2393 331
rect 2390 292 2393 328
rect 2422 302 2425 338
rect 2438 332 2441 338
rect 2446 332 2449 348
rect 2470 342 2473 398
rect 2494 392 2497 448
rect 2510 421 2513 498
rect 2518 492 2521 528
rect 2526 492 2529 518
rect 2558 482 2561 488
rect 2506 418 2513 421
rect 2530 448 2534 451
rect 2478 372 2481 378
rect 2502 342 2505 418
rect 2518 352 2521 448
rect 2536 403 2538 407
rect 2542 403 2545 407
rect 2549 403 2552 407
rect 2510 342 2513 348
rect 2462 332 2465 338
rect 2490 328 2494 331
rect 2470 292 2473 308
rect 2486 292 2489 318
rect 2502 302 2505 338
rect 2526 292 2529 358
rect 2550 352 2553 358
rect 2358 262 2361 288
rect 2518 282 2521 288
rect 2434 278 2438 281
rect 2382 262 2385 278
rect 2534 272 2537 338
rect 2490 268 2494 271
rect 2506 268 2510 271
rect 2526 268 2534 271
rect 2406 262 2409 268
rect 2450 258 2454 261
rect 2350 212 2353 258
rect 2398 252 2401 258
rect 2470 252 2473 268
rect 2478 252 2481 258
rect 2434 248 2438 251
rect 2374 181 2377 218
rect 2382 192 2385 208
rect 2374 178 2382 181
rect 2354 158 2358 161
rect 2302 152 2305 158
rect 2298 148 2302 151
rect 2362 148 2366 151
rect 2082 138 2086 141
rect 2162 138 2166 141
rect 1978 118 1982 121
rect 1962 78 1969 81
rect 1966 72 1969 78
rect 1974 62 1977 98
rect 1982 72 1985 78
rect 1998 62 2001 138
rect 2006 82 2009 118
rect 2024 103 2026 107
rect 2030 103 2033 107
rect 2037 103 2040 107
rect 2046 91 2049 98
rect 2042 88 2049 91
rect 2018 78 2022 81
rect 2030 72 2033 78
rect 2046 72 2049 78
rect 2054 62 2057 138
rect 2070 132 2073 138
rect 2150 132 2153 138
rect 2206 132 2209 138
rect 2230 132 2233 138
rect 2106 128 2110 131
rect 2138 128 2142 131
rect 2170 128 2174 131
rect 2182 122 2185 128
rect 2094 92 2097 108
rect 2062 72 2065 78
rect 2110 72 2113 118
rect 2190 92 2193 108
rect 2254 92 2257 108
rect 2270 92 2273 138
rect 2294 131 2297 138
rect 2286 128 2297 131
rect 2286 102 2289 128
rect 2294 92 2297 98
rect 2326 92 2329 148
rect 2334 112 2337 148
rect 2374 112 2377 168
rect 2390 162 2393 208
rect 2398 152 2401 238
rect 2422 152 2425 218
rect 2470 192 2473 238
rect 2510 222 2513 258
rect 2518 192 2521 268
rect 2526 202 2529 268
rect 2542 262 2545 298
rect 2550 222 2553 348
rect 2558 332 2561 338
rect 2558 242 2561 328
rect 2566 272 2569 478
rect 2582 472 2585 538
rect 2590 512 2593 538
rect 2606 532 2609 548
rect 2606 492 2609 528
rect 2614 512 2617 548
rect 2622 472 2625 538
rect 2630 532 2633 538
rect 2638 521 2641 558
rect 2646 552 2649 558
rect 2686 552 2689 558
rect 2674 548 2678 551
rect 2714 548 2718 551
rect 2678 522 2681 538
rect 2630 518 2641 521
rect 2658 518 2662 521
rect 2630 492 2633 518
rect 2662 492 2665 498
rect 2654 482 2657 488
rect 2662 482 2665 488
rect 2642 478 2646 481
rect 2670 472 2673 478
rect 2602 468 2606 471
rect 2574 392 2577 398
rect 2590 392 2593 428
rect 2586 348 2590 351
rect 2598 351 2601 458
rect 2606 362 2609 368
rect 2614 362 2617 458
rect 2622 422 2625 468
rect 2686 462 2689 538
rect 2694 512 2697 538
rect 2702 532 2705 548
rect 2726 532 2729 558
rect 2734 552 2737 558
rect 2742 552 2745 568
rect 2774 562 2777 638
rect 2758 552 2761 558
rect 2746 538 2750 541
rect 2702 492 2705 518
rect 2710 492 2713 528
rect 2774 502 2777 518
rect 2782 492 2785 528
rect 2790 492 2793 718
rect 2806 692 2809 708
rect 2814 672 2817 698
rect 2846 692 2849 738
rect 2854 732 2857 738
rect 2818 658 2822 661
rect 2798 592 2801 658
rect 2838 652 2841 658
rect 2846 632 2849 638
rect 2854 552 2857 698
rect 2862 672 2865 718
rect 2870 682 2873 738
rect 2966 732 2969 778
rect 2974 742 2977 748
rect 2982 712 2985 748
rect 2894 672 2897 708
rect 2958 692 2961 708
rect 2990 702 2993 848
rect 2998 842 3001 848
rect 3018 838 3022 841
rect 3054 752 3057 878
rect 3062 832 3065 1048
rect 3078 1022 3081 1128
rect 3086 1092 3089 1148
rect 3118 1141 3121 1148
rect 3150 1142 3153 1148
rect 3106 1138 3121 1141
rect 3138 1138 3142 1141
rect 3094 1132 3097 1138
rect 3110 1092 3113 1128
rect 3126 1102 3129 1138
rect 3158 1112 3161 1148
rect 3166 1122 3169 1248
rect 3174 1162 3177 1168
rect 3178 1148 3182 1151
rect 3194 1148 3198 1151
rect 3218 1138 3222 1141
rect 3182 1132 3185 1138
rect 3230 1132 3233 1148
rect 3238 1132 3241 1258
rect 3246 1152 3249 1258
rect 3202 1128 3206 1131
rect 3214 1112 3217 1128
rect 3262 1122 3265 1158
rect 3214 1092 3217 1108
rect 3238 1092 3241 1118
rect 3162 1078 3166 1081
rect 3086 1042 3089 1078
rect 3098 1058 3102 1061
rect 3074 948 3078 951
rect 3098 948 3102 951
rect 3110 942 3113 978
rect 3082 938 3086 941
rect 3074 928 3078 931
rect 3102 922 3105 928
rect 3118 922 3121 1078
rect 3150 1072 3153 1078
rect 3126 1052 3129 1058
rect 3154 1048 3158 1051
rect 3166 1051 3169 1068
rect 3174 1062 3177 1068
rect 3166 1048 3177 1051
rect 3126 941 3129 1048
rect 3174 1042 3177 1048
rect 3182 1042 3185 1068
rect 3198 1052 3201 1078
rect 3206 1052 3209 1078
rect 3246 1062 3249 1068
rect 3230 1052 3233 1058
rect 3254 1052 3257 1068
rect 3142 1022 3145 1028
rect 3134 952 3137 988
rect 3154 958 3158 961
rect 3142 942 3145 948
rect 3166 942 3169 988
rect 3174 942 3177 948
rect 3126 938 3137 941
rect 3106 918 3113 921
rect 3102 882 3105 888
rect 3070 821 3073 878
rect 3078 872 3081 878
rect 3110 862 3113 918
rect 3126 882 3129 928
rect 3134 892 3137 938
rect 3162 928 3166 931
rect 3166 892 3169 918
rect 3182 882 3185 1008
rect 3198 1002 3201 1038
rect 3230 1032 3233 1048
rect 3262 1032 3265 1058
rect 3190 962 3193 968
rect 3190 942 3193 948
rect 3198 942 3201 998
rect 3206 992 3209 1028
rect 3270 1012 3273 1258
rect 3294 1252 3297 1268
rect 3282 1248 3286 1251
rect 3294 1222 3297 1248
rect 3302 1172 3305 1318
rect 3310 1262 3313 1268
rect 3342 1262 3345 1348
rect 3350 1342 3353 1358
rect 3374 1351 3377 1428
rect 3370 1348 3377 1351
rect 3358 1331 3361 1338
rect 3354 1328 3361 1331
rect 3366 1302 3369 1348
rect 3382 1342 3385 1418
rect 3402 1388 3406 1391
rect 3374 1332 3377 1338
rect 3374 1291 3377 1298
rect 3366 1288 3377 1291
rect 3430 1292 3433 1438
rect 3454 1422 3457 1458
rect 3446 1418 3454 1421
rect 3438 1342 3441 1358
rect 3446 1312 3449 1418
rect 3462 1412 3465 1498
rect 3470 1452 3473 1478
rect 3478 1472 3481 1528
rect 3486 1492 3489 1548
rect 3494 1532 3497 1618
rect 3510 1602 3513 1648
rect 3506 1588 3510 1591
rect 3510 1572 3513 1578
rect 3506 1528 3510 1531
rect 3518 1492 3521 1628
rect 3526 1542 3529 1608
rect 3542 1562 3545 1708
rect 3550 1562 3553 1718
rect 3558 1572 3561 1718
rect 3538 1548 3542 1551
rect 3550 1538 3558 1541
rect 3506 1478 3510 1481
rect 3542 1472 3545 1478
rect 3522 1468 3526 1471
rect 3498 1458 3502 1461
rect 3454 1392 3457 1408
rect 3470 1382 3473 1448
rect 3542 1422 3545 1448
rect 3550 1442 3553 1538
rect 3558 1452 3561 1468
rect 3542 1392 3545 1408
rect 3470 1361 3473 1378
rect 3498 1368 3502 1371
rect 3526 1362 3529 1368
rect 3534 1362 3537 1378
rect 3462 1358 3473 1361
rect 3454 1342 3457 1348
rect 3462 1342 3465 1358
rect 3470 1342 3473 1348
rect 3478 1342 3481 1358
rect 3510 1352 3513 1358
rect 3534 1342 3537 1348
rect 3498 1338 3502 1341
rect 3546 1338 3550 1341
rect 3470 1332 3473 1338
rect 3490 1328 3494 1331
rect 3366 1272 3369 1288
rect 3462 1282 3465 1318
rect 3418 1278 3422 1281
rect 3374 1262 3377 1278
rect 3398 1262 3401 1268
rect 3350 1252 3353 1258
rect 3358 1252 3361 1258
rect 3374 1252 3377 1258
rect 3394 1248 3398 1251
rect 3342 1232 3345 1238
rect 3326 1222 3329 1228
rect 3350 1161 3353 1218
rect 3406 1192 3409 1278
rect 3478 1272 3481 1288
rect 3558 1272 3561 1288
rect 3418 1268 3422 1271
rect 3446 1262 3449 1268
rect 3434 1258 3438 1261
rect 3398 1172 3401 1178
rect 3446 1172 3449 1218
rect 3406 1162 3409 1168
rect 3350 1158 3361 1161
rect 3346 1148 3350 1151
rect 3326 1142 3329 1148
rect 3358 1142 3361 1158
rect 3366 1152 3369 1158
rect 3374 1142 3377 1158
rect 3406 1152 3409 1158
rect 3382 1142 3385 1148
rect 3346 1138 3350 1141
rect 3278 1052 3281 1108
rect 3294 1092 3297 1098
rect 3286 1082 3289 1088
rect 3302 1072 3305 1118
rect 3286 1062 3289 1068
rect 3310 1062 3313 1098
rect 3318 1062 3321 1138
rect 3338 1078 3342 1081
rect 3326 1062 3329 1068
rect 3318 1042 3321 1058
rect 3338 1048 3342 1051
rect 3350 1042 3353 1068
rect 3382 1062 3385 1088
rect 3414 1072 3417 1158
rect 3462 1151 3465 1158
rect 3430 1132 3433 1148
rect 3478 1142 3481 1268
rect 3494 1252 3497 1259
rect 3558 1172 3561 1178
rect 3526 1152 3529 1168
rect 3530 1148 3534 1151
rect 3430 1082 3433 1088
rect 3478 1072 3481 1138
rect 3410 1058 3414 1061
rect 3358 1052 3361 1058
rect 3398 1052 3401 1058
rect 3462 1052 3465 1059
rect 3370 1048 3374 1051
rect 3350 1031 3353 1038
rect 3350 1028 3361 1031
rect 3210 948 3214 951
rect 3242 948 3246 951
rect 3230 942 3233 948
rect 3278 942 3281 947
rect 3218 938 3222 941
rect 3242 938 3246 941
rect 3246 892 3249 928
rect 3254 892 3257 908
rect 3302 892 3305 968
rect 3342 962 3345 968
rect 3350 952 3353 968
rect 3310 942 3313 948
rect 3350 932 3353 938
rect 3358 892 3361 1028
rect 3406 992 3409 1038
rect 3394 968 3398 971
rect 3366 958 3393 961
rect 3366 952 3369 958
rect 3390 952 3393 958
rect 3406 952 3409 968
rect 3374 932 3377 938
rect 3382 922 3385 948
rect 3406 932 3409 948
rect 3162 878 3166 881
rect 3086 852 3089 858
rect 3126 852 3129 878
rect 3206 871 3209 888
rect 3218 878 3222 881
rect 3278 872 3281 878
rect 3334 872 3337 878
rect 3342 872 3345 888
rect 3390 882 3393 908
rect 3406 892 3409 918
rect 3390 872 3393 878
rect 3206 868 3214 871
rect 3286 862 3289 868
rect 3342 862 3345 868
rect 3174 852 3177 858
rect 3230 852 3233 858
rect 3062 818 3073 821
rect 3062 792 3065 818
rect 3078 762 3081 808
rect 3126 792 3129 838
rect 3134 802 3137 848
rect 3254 822 3257 848
rect 3398 802 3401 868
rect 3414 862 3417 1008
rect 3422 982 3425 988
rect 3462 951 3465 958
rect 3430 932 3433 948
rect 3446 921 3449 938
rect 3438 918 3449 921
rect 3438 892 3441 918
rect 3418 858 3422 861
rect 3102 772 3105 778
rect 3090 768 3094 771
rect 3034 748 3038 751
rect 3026 738 3030 741
rect 3006 732 3009 738
rect 3054 732 3057 738
rect 2998 712 3001 718
rect 3014 701 3017 718
rect 3014 698 3025 701
rect 2926 682 2929 688
rect 3006 672 3009 678
rect 3014 672 3017 688
rect 3022 682 3025 698
rect 2934 668 2942 671
rect 2978 668 2982 671
rect 2862 592 2865 668
rect 2862 562 2865 578
rect 2870 572 2873 618
rect 2878 592 2881 668
rect 2890 658 2894 661
rect 2902 642 2905 658
rect 2922 648 2926 651
rect 2802 548 2806 551
rect 2810 538 2814 541
rect 2842 538 2849 541
rect 2806 522 2809 528
rect 2814 502 2817 538
rect 2734 482 2737 488
rect 2742 482 2745 488
rect 2774 482 2777 488
rect 2722 478 2726 481
rect 2766 472 2769 478
rect 2790 472 2793 478
rect 2806 472 2809 478
rect 2642 458 2646 461
rect 2690 448 2694 451
rect 2622 352 2625 418
rect 2654 392 2657 448
rect 2702 431 2705 458
rect 2746 448 2750 451
rect 2758 442 2761 458
rect 2714 438 2718 441
rect 2702 428 2713 431
rect 2678 372 2681 418
rect 2710 392 2713 428
rect 2750 392 2753 438
rect 2694 358 2702 361
rect 2678 352 2681 358
rect 2598 348 2609 351
rect 2578 338 2582 341
rect 2606 331 2609 348
rect 2638 342 2641 348
rect 2654 342 2657 348
rect 2622 332 2625 338
rect 2606 328 2614 331
rect 2574 322 2577 328
rect 2590 292 2593 298
rect 2536 203 2538 207
rect 2542 203 2545 207
rect 2549 203 2552 207
rect 2566 202 2569 258
rect 2594 248 2598 251
rect 2566 192 2569 198
rect 2438 162 2441 168
rect 2450 158 2454 161
rect 2502 152 2505 158
rect 2406 132 2409 148
rect 2590 142 2593 238
rect 2606 192 2609 328
rect 2630 302 2633 338
rect 2634 278 2638 281
rect 2670 272 2673 338
rect 2686 332 2689 338
rect 2686 282 2689 328
rect 2634 268 2638 271
rect 2614 242 2617 258
rect 2418 138 2422 141
rect 2350 92 2353 108
rect 2398 92 2401 98
rect 2126 72 2129 88
rect 2190 75 2194 78
rect 2382 78 2401 81
rect 2414 81 2417 98
rect 2410 78 2417 81
rect 2286 72 2289 78
rect 2234 68 2238 71
rect 2158 62 2161 68
rect 1858 58 1905 61
rect 2146 58 2150 61
rect 1910 52 1913 58
rect 1954 48 1958 51
rect 1870 42 1873 48
rect 1990 42 1993 58
rect 2118 52 2121 58
rect 1842 38 1846 41
rect 2206 22 2209 68
rect 2262 62 2265 68
rect 2286 62 2289 68
rect 2218 58 2222 61
rect 2234 58 2238 61
rect 2278 58 2286 61
rect 2254 52 2257 58
rect 1486 -22 1490 -18
rect 1542 -22 1546 -18
rect 1598 -22 1602 -18
rect 1782 -22 1786 -18
rect 2134 -19 2137 18
rect 2206 -18 2209 18
rect 2278 -18 2281 58
rect 2302 42 2305 78
rect 2314 68 2318 71
rect 2326 52 2329 58
rect 2334 52 2337 68
rect 2362 58 2366 61
rect 2374 52 2377 78
rect 2382 62 2385 78
rect 2398 71 2401 78
rect 2398 68 2406 71
rect 2390 62 2393 68
rect 2410 48 2414 51
rect 2362 28 2366 31
rect 2422 22 2425 128
rect 2438 82 2441 138
rect 2486 132 2489 138
rect 2498 128 2502 131
rect 2478 122 2481 128
rect 2454 102 2457 118
rect 2446 92 2449 98
rect 2510 92 2513 138
rect 2566 122 2569 135
rect 2590 92 2593 128
rect 2606 102 2609 178
rect 2614 102 2617 128
rect 2622 122 2625 268
rect 2662 262 2665 268
rect 2670 251 2673 268
rect 2662 248 2673 251
rect 2662 192 2665 248
rect 2678 242 2681 278
rect 2694 212 2697 358
rect 2710 352 2713 368
rect 2718 342 2721 368
rect 2734 292 2737 358
rect 2746 348 2750 351
rect 2750 322 2753 348
rect 2766 312 2769 468
rect 2798 442 2801 458
rect 2814 412 2817 488
rect 2830 482 2833 488
rect 2838 482 2841 498
rect 2846 462 2849 538
rect 2862 521 2865 558
rect 2870 532 2873 538
rect 2862 518 2873 521
rect 2850 458 2854 461
rect 2790 392 2793 408
rect 2830 402 2833 448
rect 2862 432 2865 478
rect 2806 378 2825 381
rect 2806 362 2809 378
rect 2814 362 2817 368
rect 2810 348 2814 351
rect 2782 342 2785 348
rect 2774 332 2777 338
rect 2822 322 2825 378
rect 2834 348 2838 351
rect 2846 342 2849 418
rect 2870 412 2873 518
rect 2878 482 2881 548
rect 2886 542 2889 638
rect 2926 622 2929 628
rect 2934 622 2937 668
rect 2950 662 2953 668
rect 2942 658 2950 661
rect 2886 472 2889 538
rect 2902 532 2905 618
rect 2926 562 2929 568
rect 2914 548 2918 551
rect 2926 542 2929 548
rect 2910 492 2913 528
rect 2934 492 2937 618
rect 2942 532 2945 658
rect 2958 632 2961 648
rect 2974 622 2977 658
rect 2990 642 2993 658
rect 2998 612 3001 668
rect 3022 612 3025 658
rect 3030 622 3033 708
rect 3040 703 3042 707
rect 3046 703 3049 707
rect 3053 703 3056 707
rect 3038 642 3041 678
rect 3046 642 3049 658
rect 2990 592 2993 598
rect 2958 552 2961 568
rect 3002 558 3006 561
rect 2966 552 2969 558
rect 2950 542 2953 548
rect 2946 528 2950 531
rect 2974 472 2977 558
rect 3014 552 3017 558
rect 2994 548 2998 551
rect 3002 548 3006 551
rect 2982 542 2985 548
rect 3010 538 3017 541
rect 2998 492 3001 508
rect 2930 468 2934 471
rect 2878 452 2881 458
rect 2886 432 2889 468
rect 2958 462 2961 468
rect 2990 462 2993 468
rect 2910 452 2913 458
rect 2898 448 2902 451
rect 2930 448 2934 451
rect 2902 392 2905 408
rect 2950 402 2953 458
rect 2966 422 2969 448
rect 2950 392 2953 398
rect 2858 368 2862 371
rect 2870 352 2873 358
rect 2958 352 2961 358
rect 2882 348 2886 351
rect 2946 348 2953 351
rect 2854 342 2857 348
rect 2838 322 2841 338
rect 2750 292 2753 308
rect 2706 278 2710 281
rect 2702 262 2705 278
rect 2734 272 2737 288
rect 2722 268 2734 271
rect 2710 242 2713 268
rect 2782 262 2785 268
rect 2790 262 2793 318
rect 2806 292 2809 318
rect 2870 292 2873 348
rect 2890 338 2894 341
rect 2906 338 2910 341
rect 2938 338 2942 341
rect 2950 332 2953 348
rect 2962 328 2966 331
rect 2894 292 2897 308
rect 2902 301 2905 328
rect 2910 312 2913 328
rect 2958 312 2961 318
rect 2982 312 2985 458
rect 2998 412 3001 448
rect 2998 342 3001 388
rect 3006 352 3009 368
rect 2990 322 2993 328
rect 2918 301 2921 308
rect 2902 298 2921 301
rect 2818 278 2822 281
rect 2802 268 2806 271
rect 2814 261 2817 268
rect 2810 258 2817 261
rect 2726 252 2729 258
rect 2694 192 2697 208
rect 2710 162 2713 238
rect 2718 222 2721 228
rect 2666 158 2670 161
rect 2646 132 2649 138
rect 2654 122 2657 148
rect 2458 78 2462 81
rect 2502 78 2505 88
rect 2566 82 2569 88
rect 2438 62 2441 68
rect 2454 62 2457 78
rect 2478 72 2481 78
rect 2554 68 2558 71
rect 2466 58 2470 61
rect 2430 52 2433 58
rect 2334 -18 2337 8
rect 2366 -18 2369 8
rect 2414 -18 2417 8
rect 2478 -18 2481 68
rect 2546 58 2550 61
rect 2550 52 2553 58
rect 2566 22 2569 78
rect 2594 68 2598 71
rect 2606 62 2609 98
rect 2614 82 2617 98
rect 2630 82 2633 88
rect 2654 72 2657 118
rect 2646 62 2649 68
rect 2662 62 2665 108
rect 2670 102 2673 138
rect 2694 132 2698 135
rect 2678 92 2681 98
rect 2690 78 2694 81
rect 2718 72 2721 88
rect 2726 72 2729 188
rect 2734 132 2737 158
rect 2742 92 2745 198
rect 2750 152 2753 258
rect 2822 252 2825 258
rect 2774 192 2777 218
rect 2758 162 2761 178
rect 2790 162 2793 248
rect 2846 202 2849 268
rect 2854 262 2857 268
rect 2870 262 2873 288
rect 2878 272 2881 288
rect 2918 282 2921 288
rect 2974 282 2977 288
rect 2930 278 2934 281
rect 2950 272 2953 278
rect 2906 268 2910 271
rect 2930 268 2934 271
rect 2870 232 2873 248
rect 2842 158 2846 161
rect 2838 152 2841 158
rect 2862 152 2865 228
rect 2878 161 2881 268
rect 2890 258 2894 261
rect 2886 192 2889 228
rect 2926 182 2929 268
rect 2938 258 2942 261
rect 2954 248 2958 251
rect 2942 192 2945 238
rect 2966 211 2969 278
rect 2990 272 2993 298
rect 3006 292 3009 348
rect 3014 292 3017 538
rect 3022 482 3025 608
rect 3046 562 3049 618
rect 3054 602 3057 648
rect 3062 582 3065 748
rect 3078 682 3081 758
rect 3102 752 3105 758
rect 3110 712 3113 758
rect 3118 742 3121 758
rect 3142 752 3145 768
rect 3182 762 3185 768
rect 3214 762 3217 778
rect 3162 758 3166 761
rect 3214 752 3217 758
rect 3186 748 3190 751
rect 3226 748 3230 751
rect 3262 751 3265 768
rect 3290 748 3294 751
rect 3194 738 3198 741
rect 3230 732 3233 738
rect 3158 712 3161 728
rect 3110 692 3113 708
rect 3142 692 3145 708
rect 3174 692 3177 728
rect 3198 722 3201 728
rect 3198 692 3201 708
rect 3206 702 3209 718
rect 3106 678 3110 681
rect 3082 668 3086 671
rect 3074 658 3078 661
rect 3094 581 3097 678
rect 3150 672 3153 678
rect 3110 662 3113 668
rect 3118 662 3121 668
rect 3158 662 3161 688
rect 3166 662 3169 668
rect 3182 662 3185 668
rect 3130 658 3134 661
rect 3210 658 3214 661
rect 3118 651 3121 658
rect 3118 648 3129 651
rect 3102 632 3105 638
rect 3110 592 3113 598
rect 3094 578 3105 581
rect 3090 568 3094 571
rect 3102 562 3105 578
rect 3114 568 3118 571
rect 3058 558 3065 561
rect 3030 552 3033 558
rect 3034 538 3038 541
rect 3040 503 3042 507
rect 3046 503 3049 507
rect 3053 503 3056 507
rect 3038 472 3041 478
rect 3030 392 3033 438
rect 3026 368 3030 371
rect 3030 342 3033 348
rect 3046 342 3049 358
rect 3022 338 3030 341
rect 2998 262 3001 268
rect 2962 208 2969 211
rect 2870 158 2881 161
rect 2906 158 2910 161
rect 2922 158 2929 161
rect 2938 158 2942 161
rect 2766 148 2774 151
rect 2850 148 2854 151
rect 2750 132 2753 138
rect 2766 122 2769 148
rect 2806 142 2809 148
rect 2830 142 2833 148
rect 2870 142 2873 158
rect 2926 152 2929 158
rect 2882 148 2886 151
rect 2778 138 2782 141
rect 2882 138 2886 141
rect 2906 138 2910 141
rect 2810 128 2814 131
rect 2826 128 2830 131
rect 2774 92 2777 108
rect 2750 72 2753 78
rect 2758 72 2761 88
rect 2674 68 2678 71
rect 2774 62 2777 68
rect 2666 58 2670 61
rect 2698 58 2702 61
rect 2714 58 2718 61
rect 2730 58 2734 61
rect 2790 61 2793 118
rect 2894 92 2897 108
rect 2918 82 2921 148
rect 2950 142 2953 168
rect 2958 142 2961 208
rect 2982 191 2985 258
rect 3006 192 3009 268
rect 3022 262 3025 338
rect 3054 322 3057 458
rect 3062 422 3065 558
rect 3070 511 3073 548
rect 3082 538 3086 541
rect 3094 522 3097 528
rect 3070 508 3081 511
rect 3070 472 3073 488
rect 3078 442 3081 508
rect 3094 472 3097 488
rect 3102 472 3105 558
rect 3110 482 3113 518
rect 3118 492 3121 548
rect 3110 472 3113 478
rect 3114 458 3118 461
rect 3086 452 3089 458
rect 3114 448 3118 451
rect 3126 432 3129 648
rect 3134 642 3137 648
rect 3190 642 3193 658
rect 3222 652 3225 668
rect 3258 659 3262 662
rect 3286 662 3289 748
rect 3326 722 3329 728
rect 3314 688 3318 691
rect 3318 662 3321 688
rect 3334 682 3337 708
rect 3358 702 3361 747
rect 3366 672 3369 678
rect 3330 668 3334 671
rect 3210 638 3214 641
rect 3342 622 3345 658
rect 3282 588 3286 591
rect 3138 568 3142 571
rect 3242 558 3246 561
rect 3162 548 3166 551
rect 3194 548 3198 551
rect 3282 548 3286 551
rect 3322 548 3326 551
rect 3182 542 3185 548
rect 3150 502 3153 538
rect 3190 532 3193 538
rect 3222 532 3225 538
rect 3166 472 3169 528
rect 3182 522 3185 528
rect 3190 492 3193 528
rect 3214 522 3217 528
rect 3202 518 3206 521
rect 3198 492 3201 508
rect 3230 502 3233 548
rect 3342 542 3345 548
rect 3290 538 3294 541
rect 3302 531 3305 538
rect 3294 528 3305 531
rect 3326 532 3329 538
rect 3342 532 3345 538
rect 3246 522 3249 528
rect 3222 482 3225 488
rect 3250 478 3254 481
rect 3278 472 3281 498
rect 3294 472 3297 528
rect 3350 492 3353 668
rect 3374 662 3377 798
rect 3390 742 3393 748
rect 3406 662 3409 858
rect 3422 792 3425 848
rect 3438 752 3441 818
rect 3470 792 3473 808
rect 3478 782 3481 1068
rect 3494 872 3497 1098
rect 3522 1088 3526 1091
rect 3558 1042 3561 1048
rect 3526 992 3529 998
rect 3558 992 3561 998
rect 3530 948 3534 951
rect 3510 861 3513 928
rect 3522 868 3526 871
rect 3506 858 3513 861
rect 3526 852 3529 858
rect 3558 842 3561 848
rect 3494 792 3497 828
rect 3554 788 3558 791
rect 3478 752 3481 758
rect 3502 752 3505 788
rect 3518 782 3521 788
rect 3430 732 3433 748
rect 3422 712 3425 718
rect 3422 682 3425 688
rect 3438 672 3441 748
rect 3446 742 3449 748
rect 3454 722 3457 748
rect 3526 692 3529 748
rect 3514 688 3518 691
rect 3418 668 3422 671
rect 3358 652 3361 658
rect 3366 592 3369 638
rect 3390 562 3393 618
rect 3406 592 3409 658
rect 3374 532 3377 538
rect 3338 478 3342 481
rect 3146 468 3150 471
rect 3234 468 3238 471
rect 3314 468 3321 471
rect 3330 468 3334 471
rect 3142 432 3145 458
rect 3082 428 3086 431
rect 3086 412 3089 418
rect 3078 352 3081 408
rect 3066 348 3070 351
rect 3086 342 3089 408
rect 3106 368 3110 371
rect 3122 348 3126 351
rect 3070 332 3073 338
rect 3062 328 3070 331
rect 3040 303 3042 307
rect 3046 303 3049 307
rect 3053 303 3056 307
rect 3062 282 3065 328
rect 3070 292 3073 318
rect 3094 292 3097 348
rect 3134 342 3137 428
rect 3158 422 3161 468
rect 3166 452 3169 468
rect 3146 388 3150 391
rect 3166 381 3169 448
rect 3174 432 3177 458
rect 3190 422 3193 448
rect 3178 388 3182 391
rect 3166 378 3177 381
rect 3158 362 3161 368
rect 3162 348 3166 351
rect 3122 338 3126 341
rect 3102 322 3105 328
rect 3142 312 3145 348
rect 3166 312 3169 338
rect 3174 302 3177 378
rect 3198 372 3201 448
rect 3190 362 3193 368
rect 3190 352 3193 358
rect 3206 352 3209 468
rect 3246 392 3249 458
rect 3262 442 3265 458
rect 3270 392 3273 468
rect 3278 462 3281 468
rect 3322 458 3326 461
rect 3302 452 3305 458
rect 3278 392 3281 448
rect 3286 442 3289 448
rect 3246 362 3249 378
rect 3198 322 3201 338
rect 3178 278 3182 281
rect 3078 272 3081 278
rect 3126 272 3129 278
rect 3142 272 3145 278
rect 3206 272 3209 348
rect 3214 342 3217 348
rect 3222 332 3225 358
rect 3234 338 3238 341
rect 3270 341 3273 358
rect 3286 352 3289 378
rect 3266 338 3273 341
rect 3246 332 3249 338
rect 3262 332 3265 338
rect 3286 332 3289 338
rect 3294 332 3297 418
rect 3302 392 3305 448
rect 3318 352 3321 358
rect 3310 348 3318 351
rect 3310 332 3313 348
rect 3334 342 3337 428
rect 3342 422 3345 478
rect 3366 462 3369 468
rect 3374 462 3377 468
rect 3382 452 3385 518
rect 3390 492 3393 558
rect 3422 551 3425 558
rect 3438 542 3441 668
rect 3454 652 3457 659
rect 3522 658 3526 661
rect 3486 542 3489 568
rect 3494 542 3497 548
rect 3510 542 3513 548
rect 3390 461 3393 488
rect 3410 478 3414 481
rect 3454 472 3457 538
rect 3518 532 3521 548
rect 3390 458 3398 461
rect 3366 392 3369 448
rect 3398 442 3401 448
rect 3406 372 3409 378
rect 3382 352 3385 358
rect 3346 348 3350 351
rect 3374 342 3377 348
rect 3414 342 3417 348
rect 3402 338 3406 341
rect 3318 332 3321 338
rect 3222 292 3225 328
rect 3238 272 3241 278
rect 3254 272 3257 318
rect 3262 272 3265 278
rect 3162 268 3166 271
rect 3062 252 3065 258
rect 3078 242 3081 268
rect 3098 248 3102 251
rect 3022 222 3025 228
rect 3022 192 3025 218
rect 2978 188 2985 191
rect 2974 162 2977 188
rect 2990 151 2993 188
rect 3046 162 3049 188
rect 3110 172 3113 268
rect 3238 262 3241 268
rect 3126 252 3129 258
rect 3166 252 3169 258
rect 3150 242 3153 248
rect 3186 168 3190 171
rect 2986 148 2993 151
rect 3022 158 3030 161
rect 3066 158 3070 161
rect 3022 152 3025 158
rect 3034 148 3038 151
rect 3050 148 3054 151
rect 3098 148 3102 151
rect 2986 138 2990 141
rect 3090 138 3094 141
rect 2970 118 2974 121
rect 3006 92 3009 98
rect 3014 92 3017 138
rect 3022 132 3025 138
rect 3110 132 3113 138
rect 3118 132 3121 158
rect 3142 152 3145 158
rect 3130 148 3137 151
rect 3040 103 3042 107
rect 3046 103 3049 107
rect 3053 103 3056 107
rect 3062 82 3065 98
rect 3094 92 3097 98
rect 3134 92 3137 148
rect 3150 132 3153 168
rect 3198 162 3201 258
rect 3214 252 3217 258
rect 3218 248 3222 251
rect 3222 172 3225 228
rect 3162 158 3166 161
rect 3210 158 3214 161
rect 3178 148 3182 151
rect 3222 142 3225 168
rect 3158 122 3161 128
rect 3174 112 3177 138
rect 3134 82 3137 88
rect 3150 82 3153 108
rect 3182 92 3185 138
rect 3230 132 3233 178
rect 2802 78 2806 81
rect 2862 72 2865 78
rect 2942 72 2945 78
rect 3030 72 3033 78
rect 3038 72 3041 78
rect 2802 68 2806 71
rect 2930 68 2934 71
rect 2786 58 2793 61
rect 2598 52 2601 58
rect 2774 52 2777 58
rect 2586 48 2590 51
rect 2618 48 2622 51
rect 2838 42 2841 48
rect 2606 32 2609 38
rect 2854 22 2857 68
rect 2862 42 2865 68
rect 2536 3 2538 7
rect 2542 3 2545 7
rect 2549 3 2552 7
rect 2582 -18 2585 18
rect 2678 -18 2681 18
rect 2702 -18 2705 8
rect 2766 -18 2769 8
rect 2862 -18 2865 8
rect 2886 -18 2889 38
rect 2910 12 2913 68
rect 2950 62 2953 68
rect 2966 62 2969 68
rect 2918 32 2921 58
rect 2974 52 2977 68
rect 2950 42 2953 48
rect 2966 32 2969 38
rect 2982 22 2985 68
rect 3046 52 3049 78
rect 3190 75 3193 88
rect 3206 82 3209 118
rect 3222 92 3225 118
rect 3238 72 3241 208
rect 3270 192 3273 298
rect 3278 252 3281 278
rect 3294 262 3297 328
rect 3306 318 3310 321
rect 3334 291 3337 338
rect 3326 288 3337 291
rect 3350 332 3353 338
rect 3326 272 3329 288
rect 3350 278 3353 328
rect 3358 322 3361 328
rect 3358 292 3361 298
rect 3342 275 3346 278
rect 3318 252 3321 258
rect 3382 252 3385 338
rect 3422 332 3425 418
rect 3430 352 3433 468
rect 3438 382 3441 458
rect 3470 452 3473 459
rect 3506 388 3510 391
rect 3486 372 3489 378
rect 3510 352 3513 358
rect 3466 348 3470 351
rect 3438 332 3441 338
rect 3390 272 3393 308
rect 3446 302 3449 348
rect 3518 341 3521 348
rect 3514 338 3521 341
rect 3470 302 3473 328
rect 3414 272 3417 278
rect 3434 268 3438 271
rect 3246 152 3249 158
rect 3270 92 3273 178
rect 3294 152 3297 168
rect 3302 162 3305 218
rect 3342 162 3345 218
rect 3382 192 3385 248
rect 3398 242 3401 258
rect 3394 168 3398 171
rect 3278 132 3281 148
rect 3286 132 3289 148
rect 3318 132 3321 158
rect 3406 152 3409 268
rect 3414 222 3417 268
rect 3454 262 3457 268
rect 3426 258 3430 261
rect 3414 182 3417 188
rect 3422 152 3425 238
rect 3430 162 3433 168
rect 3462 152 3465 218
rect 3470 202 3473 268
rect 3494 262 3497 328
rect 3510 292 3513 338
rect 3490 258 3494 261
rect 3506 248 3510 251
rect 3478 152 3481 248
rect 3490 238 3494 241
rect 3518 192 3521 268
rect 3526 192 3529 638
rect 3538 568 3542 571
rect 3534 492 3537 528
rect 3542 512 3545 538
rect 3550 492 3553 768
rect 3558 642 3561 648
rect 3538 468 3542 471
rect 3538 348 3542 351
rect 3542 292 3545 328
rect 3542 282 3545 288
rect 3558 262 3561 518
rect 3558 252 3561 258
rect 3378 148 3382 151
rect 3342 142 3345 148
rect 3542 142 3545 208
rect 3550 152 3553 158
rect 3362 138 3366 141
rect 3482 138 3486 141
rect 3326 132 3329 138
rect 3382 132 3385 138
rect 3422 132 3425 138
rect 3454 132 3457 138
rect 3346 128 3350 131
rect 3358 128 3366 131
rect 3286 72 3289 78
rect 3130 68 3134 71
rect 3210 68 3214 71
rect 3078 42 3081 68
rect 3134 52 3137 58
rect 2910 -18 2913 8
rect 3006 -18 3009 18
rect 3150 -18 3153 68
rect 3158 42 3161 68
rect 3230 52 3233 68
rect 3294 62 3297 128
rect 3310 102 3313 118
rect 3334 112 3337 118
rect 3318 92 3321 98
rect 3358 92 3361 128
rect 3342 72 3345 78
rect 3374 72 3377 108
rect 3430 102 3433 118
rect 3462 102 3465 128
rect 3486 122 3489 128
rect 3510 102 3513 138
rect 3522 128 3526 131
rect 3462 82 3465 88
rect 3478 72 3481 78
rect 3318 52 3321 68
rect 3334 62 3337 68
rect 3378 58 3381 61
rect 3530 58 3534 61
rect 3214 42 3217 48
rect 3310 32 3313 38
rect 3526 22 3529 48
rect 3350 -18 3353 8
rect 2142 -19 2146 -18
rect 2134 -22 2146 -19
rect 2206 -22 2210 -18
rect 2278 -22 2282 -18
rect 2334 -22 2338 -18
rect 2366 -22 2370 -18
rect 2414 -22 2418 -18
rect 2478 -22 2482 -18
rect 2582 -22 2586 -18
rect 2678 -22 2682 -18
rect 2702 -22 2706 -18
rect 2766 -22 2770 -18
rect 2862 -22 2866 -18
rect 2886 -22 2890 -18
rect 2910 -22 2914 -18
rect 3006 -22 3010 -18
rect 3150 -22 3154 -18
rect 3350 -22 3354 -18
<< m3contact >>
rect 606 3298 610 3302
rect 630 3288 634 3292
rect 110 3278 114 3282
rect 254 3278 258 3282
rect 94 3268 98 3272
rect 142 3268 146 3272
rect 6 3248 10 3252
rect 30 3248 34 3252
rect 158 3248 162 3252
rect 198 3268 202 3272
rect 318 3268 322 3272
rect 222 3258 226 3262
rect 206 3248 210 3252
rect 214 3238 218 3242
rect 174 3228 178 3232
rect 102 3218 106 3222
rect 126 3218 130 3222
rect 134 3218 138 3222
rect 174 3218 178 3222
rect 78 3168 82 3172
rect 86 3168 90 3172
rect 38 3158 42 3162
rect 46 3158 50 3162
rect 118 3158 122 3162
rect 14 3138 18 3142
rect 30 3148 34 3152
rect 38 3138 42 3142
rect 22 3128 26 3132
rect 94 3148 98 3152
rect 134 3148 138 3152
rect 182 3148 186 3152
rect 86 3138 90 3142
rect 134 3138 138 3142
rect 150 3138 154 3142
rect 54 3118 58 3122
rect 158 3128 162 3132
rect 118 3118 122 3122
rect 142 3118 146 3122
rect 166 3118 170 3122
rect 174 3118 178 3122
rect 54 3088 58 3092
rect 78 3088 82 3092
rect 38 3078 42 3082
rect 62 3078 66 3082
rect 134 3078 138 3082
rect 6 3068 10 3072
rect 38 3068 42 3072
rect 78 3068 82 3072
rect 30 3058 34 3062
rect 6 3048 10 3052
rect 78 3048 82 3052
rect 22 2958 26 2962
rect 38 2948 42 2952
rect 174 3068 178 3072
rect 142 3058 146 3062
rect 86 3038 90 3042
rect 118 3038 122 3042
rect 102 2968 106 2972
rect 86 2958 90 2962
rect 134 2958 138 2962
rect 62 2948 66 2952
rect 46 2938 50 2942
rect 86 2938 90 2942
rect 38 2928 42 2932
rect 54 2928 58 2932
rect 78 2928 82 2932
rect 102 2928 106 2932
rect 22 2918 26 2922
rect 6 2878 10 2882
rect 22 2868 26 2872
rect 54 2918 58 2922
rect 198 3138 202 3142
rect 270 3258 274 3262
rect 334 3258 338 3262
rect 350 3258 354 3262
rect 366 3258 370 3262
rect 454 3268 458 3272
rect 430 3258 434 3262
rect 326 3228 330 3232
rect 318 3168 322 3172
rect 294 3148 298 3152
rect 318 3148 322 3152
rect 278 3128 282 3132
rect 294 3128 298 3132
rect 222 3118 226 3122
rect 310 3118 314 3122
rect 286 3088 290 3092
rect 190 3068 194 3072
rect 206 3068 210 3072
rect 238 3068 242 3072
rect 198 3058 202 3062
rect 206 3058 210 3062
rect 342 3248 346 3252
rect 358 3238 362 3242
rect 422 3248 426 3252
rect 478 3268 482 3272
rect 606 3268 610 3272
rect 622 3248 626 3252
rect 470 3238 474 3242
rect 518 3238 522 3242
rect 550 3238 554 3242
rect 638 3238 642 3242
rect 462 3218 466 3222
rect 398 3188 402 3192
rect 342 3168 346 3172
rect 334 3158 338 3162
rect 326 3128 330 3132
rect 318 3078 322 3082
rect 366 3128 370 3132
rect 382 3128 386 3132
rect 358 3088 362 3092
rect 350 3078 354 3082
rect 246 3058 250 3062
rect 342 3058 346 3062
rect 198 3048 202 3052
rect 222 3048 226 3052
rect 254 3048 258 3052
rect 286 3048 290 3052
rect 334 3048 338 3052
rect 270 3038 274 3042
rect 206 3028 210 3032
rect 238 3028 242 3032
rect 182 2958 186 2962
rect 190 2958 194 2962
rect 150 2948 154 2952
rect 414 3138 418 3142
rect 482 3203 486 3207
rect 489 3203 493 3207
rect 494 3188 498 3192
rect 502 3148 506 3152
rect 542 3148 546 3152
rect 462 3128 466 3132
rect 446 3118 450 3122
rect 526 3138 530 3142
rect 470 3078 474 3082
rect 398 3068 402 3072
rect 478 3068 482 3072
rect 358 3038 362 3042
rect 254 2958 258 2962
rect 278 2958 282 2962
rect 286 2958 290 2962
rect 374 2958 378 2962
rect 390 2958 394 2962
rect 238 2948 242 2952
rect 270 2948 274 2952
rect 206 2938 210 2942
rect 230 2938 234 2942
rect 174 2928 178 2932
rect 134 2918 138 2922
rect 70 2888 74 2892
rect 86 2868 90 2872
rect 94 2868 98 2872
rect 38 2858 42 2862
rect 142 2908 146 2912
rect 150 2908 154 2912
rect 110 2898 114 2902
rect 158 2878 162 2882
rect 198 2928 202 2932
rect 198 2918 202 2922
rect 190 2888 194 2892
rect 230 2918 234 2922
rect 214 2898 218 2902
rect 238 2908 242 2912
rect 262 2898 266 2902
rect 278 2898 282 2902
rect 246 2878 250 2882
rect 110 2868 114 2872
rect 150 2868 154 2872
rect 174 2868 178 2872
rect 6 2848 10 2852
rect 14 2848 18 2852
rect 70 2848 74 2852
rect 102 2848 106 2852
rect 110 2848 114 2852
rect 150 2838 154 2842
rect 94 2828 98 2832
rect 134 2828 138 2832
rect 30 2808 34 2812
rect 118 2818 122 2822
rect 166 2808 170 2812
rect 134 2768 138 2772
rect 86 2758 90 2762
rect 166 2758 170 2762
rect 174 2758 178 2762
rect 238 2868 242 2872
rect 342 2948 346 2952
rect 366 2948 370 2952
rect 310 2938 314 2942
rect 334 2938 338 2942
rect 350 2938 354 2942
rect 390 2938 394 2942
rect 294 2908 298 2912
rect 302 2898 306 2902
rect 294 2888 298 2892
rect 206 2858 210 2862
rect 246 2858 250 2862
rect 206 2848 210 2852
rect 270 2848 274 2852
rect 302 2848 306 2852
rect 286 2828 290 2832
rect 278 2758 282 2762
rect 302 2758 306 2762
rect 30 2748 34 2752
rect 14 2738 18 2742
rect 22 2728 26 2732
rect 6 2698 10 2702
rect 30 2698 34 2702
rect 14 2678 18 2682
rect 54 2748 58 2752
rect 150 2748 154 2752
rect 166 2748 170 2752
rect 150 2738 154 2742
rect 54 2728 58 2732
rect 134 2728 138 2732
rect 118 2698 122 2702
rect 94 2688 98 2692
rect 30 2668 34 2672
rect 78 2668 82 2672
rect 14 2658 18 2662
rect 22 2658 26 2662
rect 38 2658 42 2662
rect 54 2658 58 2662
rect 62 2658 66 2662
rect 86 2658 90 2662
rect 30 2648 34 2652
rect 30 2628 34 2632
rect 14 2618 18 2622
rect 6 2608 10 2612
rect 6 2558 10 2562
rect 78 2648 82 2652
rect 158 2678 162 2682
rect 446 3058 450 3062
rect 462 3058 466 3062
rect 430 3048 434 3052
rect 454 3028 458 3032
rect 582 3168 586 3172
rect 638 3168 642 3172
rect 574 3158 578 3162
rect 606 3158 610 3162
rect 598 3148 602 3152
rect 638 3148 642 3152
rect 566 3138 570 3142
rect 582 3138 586 3142
rect 558 3118 562 3122
rect 574 3118 578 3122
rect 606 3138 610 3142
rect 606 3128 610 3132
rect 598 3108 602 3112
rect 566 3098 570 3102
rect 598 3088 602 3092
rect 614 3088 618 3092
rect 670 3298 674 3302
rect 694 3298 698 3302
rect 702 3298 706 3302
rect 686 3268 690 3272
rect 670 3258 674 3262
rect 654 3218 658 3222
rect 734 3298 738 3302
rect 726 3278 730 3282
rect 710 3268 714 3272
rect 694 3258 698 3262
rect 678 3208 682 3212
rect 670 3148 674 3152
rect 662 3138 666 3142
rect 646 3108 650 3112
rect 622 3078 626 3082
rect 582 3068 586 3072
rect 558 3059 562 3063
rect 470 3048 474 3052
rect 542 3048 546 3052
rect 518 3018 522 3022
rect 482 3003 486 3007
rect 489 3003 493 3007
rect 414 2978 418 2982
rect 430 2948 434 2952
rect 534 2948 538 2952
rect 406 2938 410 2942
rect 342 2928 346 2932
rect 438 2928 442 2932
rect 318 2878 322 2882
rect 414 2918 418 2922
rect 406 2898 410 2902
rect 342 2888 346 2892
rect 334 2868 338 2872
rect 350 2868 354 2872
rect 374 2868 378 2872
rect 326 2848 330 2852
rect 366 2848 370 2852
rect 374 2798 378 2802
rect 470 2938 474 2942
rect 558 2938 562 2942
rect 446 2908 450 2912
rect 478 2908 482 2912
rect 454 2898 458 2902
rect 462 2888 466 2892
rect 470 2888 474 2892
rect 422 2878 426 2882
rect 454 2878 458 2882
rect 430 2868 434 2872
rect 462 2868 466 2872
rect 390 2858 394 2862
rect 406 2848 410 2852
rect 406 2828 410 2832
rect 382 2788 386 2792
rect 390 2778 394 2782
rect 254 2748 258 2752
rect 286 2748 290 2752
rect 310 2748 314 2752
rect 326 2748 330 2752
rect 374 2748 378 2752
rect 190 2738 194 2742
rect 190 2708 194 2712
rect 206 2738 210 2742
rect 222 2738 226 2742
rect 270 2738 274 2742
rect 278 2728 282 2732
rect 278 2718 282 2722
rect 198 2698 202 2702
rect 270 2698 274 2702
rect 214 2688 218 2692
rect 206 2678 210 2682
rect 150 2668 154 2672
rect 166 2668 170 2672
rect 190 2668 194 2672
rect 206 2668 210 2672
rect 118 2648 122 2652
rect 150 2658 154 2662
rect 166 2648 170 2652
rect 190 2648 194 2652
rect 102 2628 106 2632
rect 126 2628 130 2632
rect 182 2618 186 2622
rect 94 2608 98 2612
rect 102 2598 106 2602
rect 174 2578 178 2582
rect 78 2568 82 2572
rect 126 2568 130 2572
rect 134 2568 138 2572
rect 62 2558 66 2562
rect 78 2548 82 2552
rect 134 2548 138 2552
rect 46 2538 50 2542
rect 230 2678 234 2682
rect 246 2678 250 2682
rect 262 2678 266 2682
rect 358 2728 362 2732
rect 350 2718 354 2722
rect 366 2718 370 2722
rect 342 2708 346 2712
rect 294 2698 298 2702
rect 318 2698 322 2702
rect 326 2698 330 2702
rect 398 2768 402 2772
rect 454 2848 458 2852
rect 462 2848 466 2852
rect 446 2758 450 2762
rect 486 2848 490 2852
rect 478 2828 482 2832
rect 482 2803 486 2807
rect 489 2803 493 2807
rect 438 2748 442 2752
rect 462 2748 466 2752
rect 486 2748 490 2752
rect 598 3058 602 3062
rect 590 3028 594 3032
rect 574 2928 578 2932
rect 582 2928 586 2932
rect 734 3268 738 3272
rect 742 3268 746 3272
rect 742 3238 746 3242
rect 774 3288 778 3292
rect 782 3288 786 3292
rect 994 3303 998 3307
rect 1001 3303 1005 3307
rect 1022 3298 1026 3302
rect 1054 3298 1058 3302
rect 1142 3298 1146 3302
rect 1230 3298 1234 3302
rect 894 3288 898 3292
rect 934 3288 938 3292
rect 1014 3288 1018 3292
rect 878 3278 882 3282
rect 902 3278 906 3282
rect 966 3278 970 3282
rect 1014 3278 1018 3282
rect 1022 3278 1026 3282
rect 1086 3278 1090 3282
rect 1182 3278 1186 3282
rect 774 3268 778 3272
rect 862 3268 866 3272
rect 766 3258 770 3262
rect 862 3258 866 3262
rect 790 3248 794 3252
rect 750 3228 754 3232
rect 710 3178 714 3182
rect 734 3168 738 3172
rect 718 3158 722 3162
rect 838 3178 842 3182
rect 798 3168 802 3172
rect 822 3168 826 3172
rect 830 3168 834 3172
rect 742 3158 746 3162
rect 790 3158 794 3162
rect 886 3258 890 3262
rect 910 3258 914 3262
rect 926 3258 930 3262
rect 958 3258 962 3262
rect 942 3248 946 3252
rect 870 3238 874 3242
rect 934 3238 938 3242
rect 910 3208 914 3212
rect 774 3148 778 3152
rect 806 3148 810 3152
rect 830 3148 834 3152
rect 862 3148 866 3152
rect 702 3138 706 3142
rect 766 3138 770 3142
rect 782 3138 786 3142
rect 790 3138 794 3142
rect 798 3138 802 3142
rect 702 3128 706 3132
rect 726 3128 730 3132
rect 758 3128 762 3132
rect 686 3118 690 3122
rect 718 3118 722 3122
rect 750 3108 754 3112
rect 774 3098 778 3102
rect 678 3078 682 3082
rect 614 3058 618 3062
rect 622 3048 626 3052
rect 606 3038 610 3042
rect 686 3028 690 3032
rect 670 2998 674 3002
rect 670 2968 674 2972
rect 622 2948 626 2952
rect 630 2948 634 2952
rect 670 2948 674 2952
rect 614 2938 618 2942
rect 614 2928 618 2932
rect 630 2928 634 2932
rect 550 2878 554 2882
rect 574 2878 578 2882
rect 518 2858 522 2862
rect 542 2808 546 2812
rect 598 2858 602 2862
rect 598 2848 602 2852
rect 614 2848 618 2852
rect 582 2838 586 2842
rect 558 2798 562 2802
rect 590 2798 594 2802
rect 510 2748 514 2752
rect 542 2748 546 2752
rect 558 2748 562 2752
rect 582 2748 586 2752
rect 414 2738 418 2742
rect 502 2738 506 2742
rect 534 2738 538 2742
rect 406 2688 410 2692
rect 374 2678 378 2682
rect 286 2668 290 2672
rect 326 2668 330 2672
rect 318 2658 322 2662
rect 222 2648 226 2652
rect 222 2638 226 2642
rect 294 2648 298 2652
rect 270 2628 274 2632
rect 238 2608 242 2612
rect 262 2608 266 2612
rect 230 2588 234 2592
rect 214 2578 218 2582
rect 190 2568 194 2572
rect 238 2558 242 2562
rect 166 2538 170 2542
rect 46 2528 50 2532
rect 70 2528 74 2532
rect 30 2518 34 2522
rect 70 2518 74 2522
rect 86 2518 90 2522
rect 6 2508 10 2512
rect 6 2488 10 2492
rect 38 2498 42 2502
rect 54 2498 58 2502
rect 14 2478 18 2482
rect 30 2478 34 2482
rect 14 2468 18 2472
rect 22 2458 26 2462
rect 6 2398 10 2402
rect 46 2478 50 2482
rect 54 2478 58 2482
rect 30 2378 34 2382
rect 54 2448 58 2452
rect 62 2428 66 2432
rect 38 2368 42 2372
rect 54 2368 58 2372
rect 62 2368 66 2372
rect 46 2358 50 2362
rect 30 2348 34 2352
rect 38 2338 42 2342
rect 110 2518 114 2522
rect 158 2518 162 2522
rect 166 2518 170 2522
rect 142 2508 146 2512
rect 150 2508 154 2512
rect 158 2498 162 2502
rect 134 2478 138 2482
rect 150 2478 154 2482
rect 126 2468 130 2472
rect 94 2438 98 2442
rect 94 2378 98 2382
rect 118 2448 122 2452
rect 198 2508 202 2512
rect 206 2498 210 2502
rect 182 2488 186 2492
rect 206 2488 210 2492
rect 222 2518 226 2522
rect 310 2618 314 2622
rect 302 2578 306 2582
rect 334 2578 338 2582
rect 326 2568 330 2572
rect 318 2558 322 2562
rect 278 2548 282 2552
rect 286 2538 290 2542
rect 278 2528 282 2532
rect 286 2528 290 2532
rect 270 2508 274 2512
rect 222 2498 226 2502
rect 262 2498 266 2502
rect 174 2478 178 2482
rect 198 2478 202 2482
rect 190 2468 194 2472
rect 142 2458 146 2462
rect 166 2458 170 2462
rect 150 2448 154 2452
rect 134 2438 138 2442
rect 158 2438 162 2442
rect 110 2428 114 2432
rect 134 2428 138 2432
rect 118 2368 122 2372
rect 102 2358 106 2362
rect 110 2358 114 2362
rect 126 2358 130 2362
rect 174 2368 178 2372
rect 102 2338 106 2342
rect 78 2328 82 2332
rect 62 2298 66 2302
rect 102 2298 106 2302
rect 102 2278 106 2282
rect 126 2288 130 2292
rect 54 2268 58 2272
rect 94 2268 98 2272
rect 118 2268 122 2272
rect 22 2258 26 2262
rect 38 2258 42 2262
rect 30 2248 34 2252
rect 94 2248 98 2252
rect 54 2238 58 2242
rect 14 2168 18 2172
rect 14 2148 18 2152
rect 30 2158 34 2162
rect 78 2198 82 2202
rect 110 2178 114 2182
rect 174 2318 178 2322
rect 150 2308 154 2312
rect 150 2288 154 2292
rect 134 2268 138 2272
rect 206 2458 210 2462
rect 230 2438 234 2442
rect 238 2438 242 2442
rect 390 2678 394 2682
rect 486 2728 490 2732
rect 414 2678 418 2682
rect 414 2668 418 2672
rect 382 2658 386 2662
rect 406 2638 410 2642
rect 358 2598 362 2602
rect 358 2578 362 2582
rect 398 2598 402 2602
rect 390 2568 394 2572
rect 382 2548 386 2552
rect 470 2708 474 2712
rect 510 2708 514 2712
rect 510 2698 514 2702
rect 518 2698 522 2702
rect 446 2678 450 2682
rect 462 2678 466 2682
rect 526 2678 530 2682
rect 438 2658 442 2662
rect 446 2648 450 2652
rect 422 2608 426 2612
rect 446 2568 450 2572
rect 478 2648 482 2652
rect 462 2628 466 2632
rect 482 2603 486 2607
rect 489 2603 493 2607
rect 526 2658 530 2662
rect 518 2608 522 2612
rect 510 2578 514 2582
rect 510 2558 514 2562
rect 430 2548 434 2552
rect 470 2548 474 2552
rect 350 2538 354 2542
rect 366 2538 370 2542
rect 374 2538 378 2542
rect 326 2518 330 2522
rect 334 2518 338 2522
rect 302 2508 306 2512
rect 342 2498 346 2502
rect 326 2478 330 2482
rect 294 2468 298 2472
rect 286 2458 290 2462
rect 254 2428 258 2432
rect 238 2378 242 2382
rect 214 2358 218 2362
rect 190 2328 194 2332
rect 198 2318 202 2322
rect 222 2318 226 2322
rect 230 2318 234 2322
rect 182 2268 186 2272
rect 222 2298 226 2302
rect 134 2248 138 2252
rect 182 2248 186 2252
rect 230 2248 234 2252
rect 150 2218 154 2222
rect 166 2208 170 2212
rect 190 2168 194 2172
rect 110 2158 114 2162
rect 198 2158 202 2162
rect 214 2178 218 2182
rect 70 2148 74 2152
rect 94 2148 98 2152
rect 118 2148 122 2152
rect 206 2148 210 2152
rect 14 2128 18 2132
rect 22 2128 26 2132
rect 14 2048 18 2052
rect 6 2038 10 2042
rect 46 2068 50 2072
rect 78 2138 82 2142
rect 150 2138 154 2142
rect 158 2138 162 2142
rect 182 2138 186 2142
rect 94 2128 98 2132
rect 86 2078 90 2082
rect 70 2068 74 2072
rect 78 2058 82 2062
rect 62 2048 66 2052
rect 94 2048 98 2052
rect 46 2038 50 2042
rect 126 2108 130 2112
rect 134 2088 138 2092
rect 158 2118 162 2122
rect 174 2128 178 2132
rect 198 2128 202 2132
rect 214 2128 218 2132
rect 166 2088 170 2092
rect 166 2078 170 2082
rect 78 2028 82 2032
rect 118 2028 122 2032
rect 38 1948 42 1952
rect 6 1938 10 1942
rect 30 1938 34 1942
rect 14 1878 18 1882
rect 6 1728 10 1732
rect 70 1958 74 1962
rect 30 1868 34 1872
rect 30 1848 34 1852
rect 46 1868 50 1872
rect 94 1988 98 1992
rect 118 1968 122 1972
rect 94 1958 98 1962
rect 86 1948 90 1952
rect 126 1948 130 1952
rect 94 1938 98 1942
rect 118 1938 122 1942
rect 94 1898 98 1902
rect 102 1888 106 1892
rect 86 1868 90 1872
rect 62 1808 66 1812
rect 94 1848 98 1852
rect 78 1838 82 1842
rect 70 1798 74 1802
rect 62 1768 66 1772
rect 70 1768 74 1772
rect 30 1758 34 1762
rect 38 1748 42 1752
rect 22 1738 26 1742
rect 62 1738 66 1742
rect 38 1728 42 1732
rect 30 1708 34 1712
rect 38 1668 42 1672
rect 14 1568 18 1572
rect 38 1548 42 1552
rect 118 1908 122 1912
rect 150 2038 154 2042
rect 198 2068 202 2072
rect 246 2278 250 2282
rect 318 2438 322 2442
rect 374 2518 378 2522
rect 534 2648 538 2652
rect 534 2588 538 2592
rect 550 2708 554 2712
rect 622 2838 626 2842
rect 622 2788 626 2792
rect 622 2768 626 2772
rect 614 2738 618 2742
rect 566 2728 570 2732
rect 558 2698 562 2702
rect 558 2678 562 2682
rect 590 2688 594 2692
rect 646 2908 650 2912
rect 654 2898 658 2902
rect 678 2938 682 2942
rect 710 3008 714 3012
rect 758 3058 762 3062
rect 734 3018 738 3022
rect 734 3008 738 3012
rect 734 2998 738 3002
rect 726 2988 730 2992
rect 718 2978 722 2982
rect 710 2958 714 2962
rect 726 2958 730 2962
rect 694 2948 698 2952
rect 686 2928 690 2932
rect 806 3128 810 3132
rect 846 3128 850 3132
rect 862 3128 866 3132
rect 814 3098 818 3102
rect 846 3098 850 3102
rect 830 3088 834 3092
rect 846 3078 850 3082
rect 806 3058 810 3062
rect 798 3038 802 3042
rect 830 3028 834 3032
rect 782 2958 786 2962
rect 742 2948 746 2952
rect 790 2938 794 2942
rect 694 2918 698 2922
rect 718 2918 722 2922
rect 758 2918 762 2922
rect 830 2998 834 3002
rect 822 2948 826 2952
rect 806 2938 810 2942
rect 862 3098 866 3102
rect 870 3088 874 3092
rect 1006 3258 1010 3262
rect 1038 3258 1042 3262
rect 1054 3258 1058 3262
rect 1078 3258 1082 3262
rect 1022 3248 1026 3252
rect 1070 3248 1074 3252
rect 1054 3238 1058 3242
rect 1070 3228 1074 3232
rect 1102 3258 1106 3262
rect 1286 3298 1290 3302
rect 1350 3298 1354 3302
rect 1270 3288 1274 3292
rect 1358 3288 1362 3292
rect 1190 3258 1194 3262
rect 1246 3258 1250 3262
rect 1326 3258 1330 3262
rect 1118 3248 1122 3252
rect 1326 3248 1330 3252
rect 1294 3238 1298 3242
rect 1094 3228 1098 3232
rect 1198 3228 1202 3232
rect 1078 3198 1082 3202
rect 1110 3198 1114 3202
rect 1014 3188 1018 3192
rect 998 3178 1002 3182
rect 966 3168 970 3172
rect 1190 3168 1194 3172
rect 1022 3158 1026 3162
rect 950 3148 954 3152
rect 958 3148 962 3152
rect 966 3128 970 3132
rect 1054 3148 1058 3152
rect 1062 3148 1066 3152
rect 1110 3148 1114 3152
rect 1158 3148 1162 3152
rect 990 3138 994 3142
rect 918 3118 922 3122
rect 942 3118 946 3122
rect 974 3118 978 3122
rect 1038 3118 1042 3122
rect 910 3108 914 3112
rect 918 3098 922 3102
rect 918 3078 922 3082
rect 918 3058 922 3062
rect 910 3008 914 3012
rect 994 3103 998 3107
rect 1001 3103 1005 3107
rect 966 3098 970 3102
rect 958 3088 962 3092
rect 966 3058 970 3062
rect 1022 3058 1026 3062
rect 950 3048 954 3052
rect 934 3018 938 3022
rect 1038 3048 1042 3052
rect 1062 3138 1066 3142
rect 1126 3138 1130 3142
rect 1166 3138 1170 3142
rect 1070 3128 1074 3132
rect 1094 3118 1098 3122
rect 1118 3118 1122 3122
rect 1134 3118 1138 3122
rect 1262 3198 1266 3202
rect 1270 3178 1274 3182
rect 1246 3168 1250 3172
rect 1206 3158 1210 3162
rect 1238 3148 1242 3152
rect 1254 3148 1258 3152
rect 1190 3138 1194 3142
rect 1182 3118 1186 3122
rect 1358 3258 1362 3262
rect 1374 3258 1378 3262
rect 1342 3168 1346 3172
rect 1366 3248 1370 3252
rect 1382 3218 1386 3222
rect 1382 3158 1386 3162
rect 1286 3148 1290 3152
rect 1310 3148 1314 3152
rect 1342 3148 1346 3152
rect 1358 3148 1362 3152
rect 1278 3138 1282 3142
rect 1374 3138 1378 3142
rect 1214 3128 1218 3132
rect 1238 3128 1242 3132
rect 1230 3098 1234 3102
rect 1158 3088 1162 3092
rect 1078 3078 1082 3082
rect 1102 3078 1106 3082
rect 1134 3078 1138 3082
rect 1142 3078 1146 3082
rect 1206 3078 1210 3082
rect 1062 3058 1066 3062
rect 1118 3058 1122 3062
rect 1142 3058 1146 3062
rect 1126 3048 1130 3052
rect 1078 3038 1082 3042
rect 1086 3038 1090 3042
rect 1294 3108 1298 3112
rect 1254 3098 1258 3102
rect 1326 3088 1330 3092
rect 1286 3078 1290 3082
rect 1366 3108 1370 3112
rect 1414 3298 1418 3302
rect 1454 3258 1458 3262
rect 1430 3238 1434 3242
rect 1398 3228 1402 3232
rect 1430 3208 1434 3212
rect 1398 3178 1402 3182
rect 1398 3168 1402 3172
rect 1486 3268 1490 3272
rect 1518 3268 1522 3272
rect 1478 3258 1482 3262
rect 1502 3258 1506 3262
rect 1470 3248 1474 3252
rect 1486 3248 1490 3252
rect 1510 3238 1514 3242
rect 1518 3238 1522 3242
rect 1478 3208 1482 3212
rect 1514 3203 1518 3207
rect 1521 3203 1525 3207
rect 1462 3188 1466 3192
rect 1510 3178 1514 3182
rect 1494 3148 1498 3152
rect 1398 3118 1402 3122
rect 1446 3138 1450 3142
rect 1462 3098 1466 3102
rect 1518 3138 1522 3142
rect 1406 3088 1410 3092
rect 1430 3088 1434 3092
rect 1526 3088 1530 3092
rect 1374 3078 1378 3082
rect 1510 3078 1514 3082
rect 1118 3038 1122 3042
rect 1222 3038 1226 3042
rect 1118 3028 1122 3032
rect 1038 3018 1042 3022
rect 1046 3018 1050 3022
rect 1094 3018 1098 3022
rect 934 2988 938 2992
rect 974 2988 978 2992
rect 918 2978 922 2982
rect 854 2968 858 2972
rect 846 2958 850 2962
rect 870 2958 874 2962
rect 854 2948 858 2952
rect 806 2928 810 2932
rect 830 2928 834 2932
rect 670 2878 674 2882
rect 686 2878 690 2882
rect 782 2878 786 2882
rect 638 2868 642 2872
rect 654 2868 658 2872
rect 726 2868 730 2872
rect 766 2868 770 2872
rect 774 2868 778 2872
rect 926 2938 930 2942
rect 894 2928 898 2932
rect 910 2928 914 2932
rect 830 2888 834 2892
rect 838 2888 842 2892
rect 854 2888 858 2892
rect 822 2878 826 2882
rect 814 2868 818 2872
rect 718 2858 722 2862
rect 790 2858 794 2862
rect 686 2848 690 2852
rect 710 2848 714 2852
rect 670 2838 674 2842
rect 654 2808 658 2812
rect 638 2798 642 2802
rect 678 2798 682 2802
rect 638 2768 642 2772
rect 662 2748 666 2752
rect 718 2828 722 2832
rect 726 2828 730 2832
rect 686 2788 690 2792
rect 782 2818 786 2822
rect 726 2808 730 2812
rect 702 2748 706 2752
rect 630 2738 634 2742
rect 694 2738 698 2742
rect 758 2738 762 2742
rect 766 2738 770 2742
rect 654 2728 658 2732
rect 718 2728 722 2732
rect 734 2728 738 2732
rect 614 2698 618 2702
rect 702 2708 706 2712
rect 726 2708 730 2712
rect 654 2698 658 2702
rect 670 2698 674 2702
rect 686 2698 690 2702
rect 638 2678 642 2682
rect 694 2678 698 2682
rect 598 2658 602 2662
rect 622 2658 626 2662
rect 654 2658 658 2662
rect 598 2648 602 2652
rect 606 2648 610 2652
rect 550 2638 554 2642
rect 582 2638 586 2642
rect 590 2628 594 2632
rect 558 2598 562 2602
rect 470 2538 474 2542
rect 486 2538 490 2542
rect 518 2538 522 2542
rect 526 2538 530 2542
rect 534 2538 538 2542
rect 566 2568 570 2572
rect 582 2568 586 2572
rect 590 2558 594 2562
rect 566 2548 570 2552
rect 878 2878 882 2882
rect 846 2858 850 2862
rect 862 2858 866 2862
rect 846 2818 850 2822
rect 870 2818 874 2822
rect 798 2798 802 2802
rect 806 2798 810 2802
rect 830 2788 834 2792
rect 790 2768 794 2772
rect 822 2768 826 2772
rect 782 2738 786 2742
rect 798 2738 802 2742
rect 814 2738 818 2742
rect 846 2758 850 2762
rect 942 2978 946 2982
rect 950 2958 954 2962
rect 1022 2958 1026 2962
rect 1086 2998 1090 3002
rect 1062 2958 1066 2962
rect 966 2938 970 2942
rect 974 2938 978 2942
rect 990 2938 994 2942
rect 1014 2938 1018 2942
rect 1046 2938 1050 2942
rect 1078 2938 1082 2942
rect 1046 2928 1050 2932
rect 1046 2918 1050 2922
rect 1022 2908 1026 2912
rect 994 2903 998 2907
rect 1001 2903 1005 2907
rect 1030 2898 1034 2902
rect 950 2888 954 2892
rect 982 2888 986 2892
rect 902 2878 906 2882
rect 934 2878 938 2882
rect 910 2868 914 2872
rect 942 2868 946 2872
rect 910 2838 914 2842
rect 926 2838 930 2842
rect 886 2778 890 2782
rect 862 2758 866 2762
rect 886 2748 890 2752
rect 838 2738 842 2742
rect 750 2678 754 2682
rect 734 2658 738 2662
rect 750 2658 754 2662
rect 758 2658 762 2662
rect 766 2658 770 2662
rect 702 2648 706 2652
rect 678 2638 682 2642
rect 686 2638 690 2642
rect 718 2628 722 2632
rect 614 2588 618 2592
rect 646 2588 650 2592
rect 622 2548 626 2552
rect 614 2538 618 2542
rect 670 2538 674 2542
rect 406 2518 410 2522
rect 446 2518 450 2522
rect 462 2518 466 2522
rect 502 2518 506 2522
rect 542 2508 546 2512
rect 406 2488 410 2492
rect 398 2468 402 2472
rect 446 2478 450 2482
rect 470 2478 474 2482
rect 494 2478 498 2482
rect 438 2468 442 2472
rect 526 2468 530 2472
rect 518 2458 522 2462
rect 374 2418 378 2422
rect 350 2408 354 2412
rect 310 2398 314 2402
rect 286 2368 290 2372
rect 302 2328 306 2332
rect 278 2278 282 2282
rect 254 2248 258 2252
rect 246 2138 250 2142
rect 270 2198 274 2202
rect 278 2168 282 2172
rect 254 2128 258 2132
rect 262 2128 266 2132
rect 238 2088 242 2092
rect 174 2028 178 2032
rect 166 1968 170 1972
rect 342 2378 346 2382
rect 398 2388 402 2392
rect 478 2448 482 2452
rect 502 2448 506 2452
rect 422 2438 426 2442
rect 414 2428 418 2432
rect 454 2418 458 2422
rect 438 2378 442 2382
rect 318 2368 322 2372
rect 358 2368 362 2372
rect 374 2368 378 2372
rect 334 2328 338 2332
rect 350 2328 354 2332
rect 350 2308 354 2312
rect 334 2278 338 2282
rect 302 2248 306 2252
rect 294 2168 298 2172
rect 342 2248 346 2252
rect 334 2238 338 2242
rect 342 2178 346 2182
rect 310 2168 314 2172
rect 310 2158 314 2162
rect 334 2148 338 2152
rect 302 2088 306 2092
rect 278 2078 282 2082
rect 310 2078 314 2082
rect 326 2108 330 2112
rect 246 2068 250 2072
rect 262 2068 266 2072
rect 278 2068 282 2072
rect 318 2068 322 2072
rect 398 2338 402 2342
rect 406 2338 410 2342
rect 422 2338 426 2342
rect 438 2338 442 2342
rect 366 2328 370 2332
rect 382 2328 386 2332
rect 414 2328 418 2332
rect 430 2328 434 2332
rect 366 2268 370 2272
rect 406 2318 410 2322
rect 390 2278 394 2282
rect 438 2308 442 2312
rect 446 2268 450 2272
rect 486 2428 490 2432
rect 502 2418 506 2422
rect 482 2403 486 2407
rect 489 2403 493 2407
rect 462 2398 466 2402
rect 462 2388 466 2392
rect 470 2338 474 2342
rect 486 2328 490 2332
rect 494 2308 498 2312
rect 494 2298 498 2302
rect 574 2508 578 2512
rect 582 2508 586 2512
rect 566 2488 570 2492
rect 606 2518 610 2522
rect 686 2608 690 2612
rect 766 2648 770 2652
rect 758 2628 762 2632
rect 750 2598 754 2602
rect 726 2568 730 2572
rect 718 2548 722 2552
rect 734 2548 738 2552
rect 806 2658 810 2662
rect 806 2638 810 2642
rect 790 2628 794 2632
rect 830 2728 834 2732
rect 910 2778 914 2782
rect 1030 2878 1034 2882
rect 1054 2878 1058 2882
rect 1070 2928 1074 2932
rect 1070 2888 1074 2892
rect 982 2868 986 2872
rect 966 2858 970 2862
rect 950 2828 954 2832
rect 990 2788 994 2792
rect 934 2768 938 2772
rect 942 2768 946 2772
rect 942 2758 946 2762
rect 1014 2758 1018 2762
rect 990 2748 994 2752
rect 870 2738 874 2742
rect 894 2738 898 2742
rect 918 2738 922 2742
rect 926 2738 930 2742
rect 838 2698 842 2702
rect 878 2698 882 2702
rect 902 2698 906 2702
rect 830 2658 834 2662
rect 822 2638 826 2642
rect 814 2618 818 2622
rect 766 2608 770 2612
rect 782 2608 786 2612
rect 790 2588 794 2592
rect 854 2638 858 2642
rect 926 2698 930 2702
rect 934 2688 938 2692
rect 950 2708 954 2712
rect 942 2668 946 2672
rect 910 2658 914 2662
rect 934 2658 938 2662
rect 878 2638 882 2642
rect 918 2638 922 2642
rect 926 2638 930 2642
rect 846 2628 850 2632
rect 870 2628 874 2632
rect 886 2628 890 2632
rect 910 2628 914 2632
rect 878 2608 882 2612
rect 830 2598 834 2602
rect 878 2598 882 2602
rect 982 2738 986 2742
rect 994 2703 998 2707
rect 1001 2703 1005 2707
rect 1062 2868 1066 2872
rect 1070 2868 1074 2872
rect 1030 2848 1034 2852
rect 1030 2828 1034 2832
rect 1094 2958 1098 2962
rect 1102 2938 1106 2942
rect 1102 2928 1106 2932
rect 1222 3018 1226 3022
rect 1230 3008 1234 3012
rect 1222 2978 1226 2982
rect 1182 2968 1186 2972
rect 1118 2958 1122 2962
rect 1142 2958 1146 2962
rect 1158 2958 1162 2962
rect 1134 2938 1138 2942
rect 1174 2938 1178 2942
rect 1158 2908 1162 2912
rect 1118 2898 1122 2902
rect 1150 2898 1154 2902
rect 1110 2888 1114 2892
rect 1094 2868 1098 2872
rect 1214 2958 1218 2962
rect 1190 2938 1194 2942
rect 1222 2938 1226 2942
rect 1246 3048 1250 3052
rect 1270 3048 1274 3052
rect 1310 3048 1314 3052
rect 1238 2988 1242 2992
rect 1254 2988 1258 2992
rect 1214 2928 1218 2932
rect 1222 2928 1226 2932
rect 1134 2888 1138 2892
rect 1166 2888 1170 2892
rect 1206 2878 1210 2882
rect 1230 2878 1234 2882
rect 1238 2878 1242 2882
rect 1142 2858 1146 2862
rect 1078 2838 1082 2842
rect 1142 2848 1146 2852
rect 1118 2818 1122 2822
rect 1110 2808 1114 2812
rect 1102 2788 1106 2792
rect 1054 2728 1058 2732
rect 1062 2718 1066 2722
rect 1046 2708 1050 2712
rect 1014 2638 1018 2642
rect 982 2618 986 2622
rect 1102 2758 1106 2762
rect 1094 2738 1098 2742
rect 1134 2808 1138 2812
rect 1134 2798 1138 2802
rect 1118 2788 1122 2792
rect 1126 2748 1130 2752
rect 1102 2728 1106 2732
rect 1086 2708 1090 2712
rect 1094 2688 1098 2692
rect 1038 2658 1042 2662
rect 1062 2658 1066 2662
rect 1054 2628 1058 2632
rect 1030 2608 1034 2612
rect 958 2588 962 2592
rect 830 2578 834 2582
rect 902 2578 906 2582
rect 782 2558 786 2562
rect 806 2558 810 2562
rect 782 2548 786 2552
rect 1078 2608 1082 2612
rect 1110 2658 1114 2662
rect 1254 2938 1258 2942
rect 1278 2938 1282 2942
rect 1262 2928 1266 2932
rect 1278 2888 1282 2892
rect 1262 2878 1266 2882
rect 1310 3028 1314 3032
rect 1310 3018 1314 3022
rect 1302 3008 1306 3012
rect 1318 2968 1322 2972
rect 1366 3048 1370 3052
rect 1342 2998 1346 3002
rect 1310 2938 1314 2942
rect 1326 2938 1330 2942
rect 1182 2868 1186 2872
rect 1286 2868 1290 2872
rect 1318 2918 1322 2922
rect 1326 2918 1330 2922
rect 1350 2968 1354 2972
rect 1374 3028 1378 3032
rect 1398 3048 1402 3052
rect 1414 3048 1418 3052
rect 1390 3018 1394 3022
rect 1366 2968 1370 2972
rect 1358 2958 1362 2962
rect 1342 2928 1346 2932
rect 1350 2928 1354 2932
rect 1430 3038 1434 3042
rect 1446 3048 1450 3052
rect 1438 3028 1442 3032
rect 1422 3018 1426 3022
rect 1478 3048 1482 3052
rect 1486 3048 1490 3052
rect 1478 3018 1482 3022
rect 1430 2998 1434 3002
rect 1470 2998 1474 3002
rect 1502 3008 1506 3012
rect 1494 2998 1498 3002
rect 1454 2978 1458 2982
rect 1470 2968 1474 2972
rect 1478 2968 1482 2972
rect 1414 2958 1418 2962
rect 1430 2958 1434 2962
rect 1446 2958 1450 2962
rect 1454 2958 1458 2962
rect 1374 2918 1378 2922
rect 1174 2858 1178 2862
rect 1302 2858 1306 2862
rect 1326 2858 1330 2862
rect 1174 2848 1178 2852
rect 1198 2848 1202 2852
rect 1222 2848 1226 2852
rect 1230 2848 1234 2852
rect 1270 2848 1274 2852
rect 1310 2848 1314 2852
rect 1422 2918 1426 2922
rect 1406 2908 1410 2912
rect 1414 2908 1418 2912
rect 1454 2928 1458 2932
rect 1438 2898 1442 2902
rect 1454 2898 1458 2902
rect 1382 2868 1386 2872
rect 1398 2868 1402 2872
rect 1430 2868 1434 2872
rect 1374 2858 1378 2862
rect 1198 2838 1202 2842
rect 1150 2798 1154 2802
rect 1270 2838 1274 2842
rect 1286 2838 1290 2842
rect 1270 2798 1274 2802
rect 1286 2788 1290 2792
rect 1302 2788 1306 2792
rect 1238 2768 1242 2772
rect 1150 2758 1154 2762
rect 1198 2758 1202 2762
rect 1214 2758 1218 2762
rect 1230 2758 1234 2762
rect 1174 2748 1178 2752
rect 1214 2748 1218 2752
rect 1142 2698 1146 2702
rect 1174 2738 1178 2742
rect 1190 2728 1194 2732
rect 1230 2708 1234 2712
rect 1222 2698 1226 2702
rect 1134 2668 1138 2672
rect 1150 2668 1154 2672
rect 1166 2668 1170 2672
rect 1174 2668 1178 2672
rect 1134 2658 1138 2662
rect 1182 2658 1186 2662
rect 1214 2658 1218 2662
rect 1254 2698 1258 2702
rect 1246 2658 1250 2662
rect 1230 2648 1234 2652
rect 1382 2848 1386 2852
rect 1390 2848 1394 2852
rect 1406 2848 1410 2852
rect 1374 2838 1378 2842
rect 1350 2808 1354 2812
rect 1358 2798 1362 2802
rect 1350 2778 1354 2782
rect 1318 2748 1322 2752
rect 1302 2738 1306 2742
rect 1310 2738 1314 2742
rect 1334 2738 1338 2742
rect 1294 2728 1298 2732
rect 1326 2728 1330 2732
rect 1342 2728 1346 2732
rect 1262 2688 1266 2692
rect 1270 2678 1274 2682
rect 1270 2668 1274 2672
rect 1278 2658 1282 2662
rect 1142 2638 1146 2642
rect 1102 2618 1106 2622
rect 1086 2588 1090 2592
rect 846 2558 850 2562
rect 878 2558 882 2562
rect 1070 2558 1074 2562
rect 1110 2558 1114 2562
rect 1214 2628 1218 2632
rect 1230 2628 1234 2632
rect 1142 2588 1146 2592
rect 1182 2588 1186 2592
rect 1174 2558 1178 2562
rect 1190 2558 1194 2562
rect 1214 2558 1218 2562
rect 918 2548 922 2552
rect 942 2548 946 2552
rect 974 2548 978 2552
rect 1022 2548 1026 2552
rect 1118 2548 1122 2552
rect 1126 2548 1130 2552
rect 710 2538 714 2542
rect 750 2538 754 2542
rect 934 2538 938 2542
rect 686 2528 690 2532
rect 702 2528 706 2532
rect 742 2528 746 2532
rect 678 2518 682 2522
rect 630 2498 634 2502
rect 598 2478 602 2482
rect 606 2478 610 2482
rect 566 2458 570 2462
rect 542 2448 546 2452
rect 566 2448 570 2452
rect 534 2438 538 2442
rect 590 2448 594 2452
rect 558 2398 562 2402
rect 582 2398 586 2402
rect 582 2378 586 2382
rect 510 2348 514 2352
rect 510 2338 514 2342
rect 534 2338 538 2342
rect 526 2328 530 2332
rect 502 2268 506 2272
rect 462 2248 466 2252
rect 390 2238 394 2242
rect 358 2208 362 2212
rect 366 2168 370 2172
rect 382 2148 386 2152
rect 366 2138 370 2142
rect 414 2138 418 2142
rect 342 2118 346 2122
rect 350 2118 354 2122
rect 342 2078 346 2082
rect 262 2038 266 2042
rect 350 2038 354 2042
rect 246 2018 250 2022
rect 214 1998 218 2002
rect 174 1958 178 1962
rect 150 1948 154 1952
rect 142 1898 146 1902
rect 142 1888 146 1892
rect 110 1778 114 1782
rect 86 1758 90 1762
rect 86 1748 90 1752
rect 110 1748 114 1752
rect 78 1738 82 1742
rect 78 1698 82 1702
rect 54 1568 58 1572
rect 22 1538 26 1542
rect 30 1538 34 1542
rect 54 1538 58 1542
rect 190 1958 194 1962
rect 206 1948 210 1952
rect 174 1938 178 1942
rect 166 1928 170 1932
rect 230 1988 234 1992
rect 238 1968 242 1972
rect 262 2008 266 2012
rect 262 1978 266 1982
rect 230 1928 234 1932
rect 214 1908 218 1912
rect 206 1878 210 1882
rect 206 1868 210 1872
rect 222 1868 226 1872
rect 174 1848 178 1852
rect 150 1838 154 1842
rect 142 1778 146 1782
rect 158 1758 162 1762
rect 118 1738 122 1742
rect 158 1738 162 1742
rect 174 1728 178 1732
rect 134 1718 138 1722
rect 150 1718 154 1722
rect 110 1678 114 1682
rect 254 1918 258 1922
rect 246 1858 250 1862
rect 222 1828 226 1832
rect 254 1788 258 1792
rect 254 1768 258 1772
rect 190 1758 194 1762
rect 238 1748 242 1752
rect 198 1738 202 1742
rect 286 1988 290 1992
rect 302 1988 306 1992
rect 294 1978 298 1982
rect 278 1948 282 1952
rect 278 1938 282 1942
rect 310 1978 314 1982
rect 270 1868 274 1872
rect 334 1948 338 1952
rect 350 1938 354 1942
rect 318 1898 322 1902
rect 302 1858 306 1862
rect 318 1858 322 1862
rect 294 1838 298 1842
rect 270 1758 274 1762
rect 294 1758 298 1762
rect 278 1738 282 1742
rect 230 1728 234 1732
rect 222 1708 226 1712
rect 238 1688 242 1692
rect 238 1678 242 1682
rect 254 1678 258 1682
rect 182 1668 186 1672
rect 222 1668 226 1672
rect 158 1658 162 1662
rect 110 1648 114 1652
rect 102 1638 106 1642
rect 214 1658 218 1662
rect 190 1648 194 1652
rect 198 1648 202 1652
rect 222 1648 226 1652
rect 166 1628 170 1632
rect 166 1618 170 1622
rect 150 1608 154 1612
rect 126 1588 130 1592
rect 94 1558 98 1562
rect 102 1558 106 1562
rect 150 1568 154 1572
rect 134 1558 138 1562
rect 158 1558 162 1562
rect 118 1548 122 1552
rect 150 1548 154 1552
rect 54 1468 58 1472
rect 62 1438 66 1442
rect 78 1488 82 1492
rect 190 1568 194 1572
rect 230 1638 234 1642
rect 206 1628 210 1632
rect 214 1578 218 1582
rect 270 1678 274 1682
rect 262 1668 266 1672
rect 262 1658 266 1662
rect 270 1608 274 1612
rect 254 1568 258 1572
rect 214 1548 218 1552
rect 198 1538 202 1542
rect 158 1528 162 1532
rect 174 1528 178 1532
rect 190 1528 194 1532
rect 166 1518 170 1522
rect 174 1478 178 1482
rect 94 1468 98 1472
rect 78 1458 82 1462
rect 94 1458 98 1462
rect 102 1448 106 1452
rect 110 1448 114 1452
rect 134 1458 138 1462
rect 126 1438 130 1442
rect 54 1368 58 1372
rect 70 1368 74 1372
rect 102 1368 106 1372
rect 110 1358 114 1362
rect 46 1348 50 1352
rect 70 1348 74 1352
rect 30 1338 34 1342
rect 14 1308 18 1312
rect 14 1278 18 1282
rect 14 1258 18 1262
rect 30 1248 34 1252
rect 62 1308 66 1312
rect 206 1478 210 1482
rect 198 1468 202 1472
rect 190 1458 194 1462
rect 150 1448 154 1452
rect 166 1448 170 1452
rect 166 1438 170 1442
rect 182 1368 186 1372
rect 142 1348 146 1352
rect 166 1348 170 1352
rect 190 1348 194 1352
rect 94 1338 98 1342
rect 126 1338 130 1342
rect 110 1328 114 1332
rect 70 1288 74 1292
rect 62 1258 66 1262
rect 86 1258 90 1262
rect 70 1228 74 1232
rect 78 1208 82 1212
rect 134 1278 138 1282
rect 62 1168 66 1172
rect 94 1168 98 1172
rect 94 1158 98 1162
rect 102 1158 106 1162
rect 30 1148 34 1152
rect 6 1128 10 1132
rect 6 1118 10 1122
rect 14 1058 18 1062
rect 46 1138 50 1142
rect 102 1148 106 1152
rect 134 1248 138 1252
rect 142 1218 146 1222
rect 134 1188 138 1192
rect 166 1288 170 1292
rect 166 1268 170 1272
rect 166 1168 170 1172
rect 262 1558 266 1562
rect 254 1498 258 1502
rect 254 1448 258 1452
rect 310 1818 314 1822
rect 286 1698 290 1702
rect 318 1718 322 1722
rect 302 1678 306 1682
rect 310 1678 314 1682
rect 334 1898 338 1902
rect 334 1718 338 1722
rect 326 1678 330 1682
rect 326 1668 330 1672
rect 382 2098 386 2102
rect 406 2128 410 2132
rect 390 2058 394 2062
rect 374 1998 378 2002
rect 374 1988 378 1992
rect 382 1948 386 1952
rect 398 1948 402 1952
rect 390 1938 394 1942
rect 406 1918 410 1922
rect 382 1898 386 1902
rect 366 1868 370 1872
rect 350 1838 354 1842
rect 358 1768 362 1772
rect 350 1758 354 1762
rect 374 1838 378 1842
rect 446 2208 450 2212
rect 430 2168 434 2172
rect 446 2148 450 2152
rect 482 2203 486 2207
rect 489 2203 493 2207
rect 478 2168 482 2172
rect 478 2118 482 2122
rect 454 2108 458 2112
rect 462 2108 466 2112
rect 454 2098 458 2102
rect 422 2078 426 2082
rect 438 2078 442 2082
rect 422 2008 426 2012
rect 422 1988 426 1992
rect 430 1988 434 1992
rect 430 1978 434 1982
rect 470 2088 474 2092
rect 446 2038 450 2042
rect 462 2028 466 2032
rect 438 1958 442 1962
rect 446 1948 450 1952
rect 414 1898 418 1902
rect 430 1898 434 1902
rect 454 1898 458 1902
rect 398 1838 402 1842
rect 390 1788 394 1792
rect 382 1768 386 1772
rect 374 1758 378 1762
rect 494 2058 498 2062
rect 518 2268 522 2272
rect 550 2348 554 2352
rect 622 2458 626 2462
rect 710 2488 714 2492
rect 662 2478 666 2482
rect 678 2458 682 2462
rect 686 2458 690 2462
rect 830 2528 834 2532
rect 798 2498 802 2502
rect 774 2488 778 2492
rect 766 2478 770 2482
rect 782 2468 786 2472
rect 862 2528 866 2532
rect 894 2528 898 2532
rect 870 2518 874 2522
rect 846 2508 850 2512
rect 758 2458 762 2462
rect 790 2458 794 2462
rect 822 2458 826 2462
rect 614 2358 618 2362
rect 598 2338 602 2342
rect 614 2328 618 2332
rect 566 2318 570 2322
rect 550 2298 554 2302
rect 542 2288 546 2292
rect 574 2278 578 2282
rect 606 2308 610 2312
rect 614 2308 618 2312
rect 598 2278 602 2282
rect 550 2268 554 2272
rect 582 2268 586 2272
rect 614 2268 618 2272
rect 526 2248 530 2252
rect 678 2418 682 2422
rect 638 2368 642 2372
rect 630 2358 634 2362
rect 710 2398 714 2402
rect 766 2448 770 2452
rect 814 2448 818 2452
rect 766 2438 770 2442
rect 694 2388 698 2392
rect 726 2388 730 2392
rect 758 2398 762 2402
rect 750 2378 754 2382
rect 702 2368 706 2372
rect 734 2368 738 2372
rect 662 2358 666 2362
rect 726 2358 730 2362
rect 758 2358 762 2362
rect 678 2348 682 2352
rect 654 2338 658 2342
rect 670 2338 674 2342
rect 686 2338 690 2342
rect 646 2318 650 2322
rect 630 2298 634 2302
rect 614 2258 618 2262
rect 574 2248 578 2252
rect 646 2248 650 2252
rect 590 2238 594 2242
rect 558 2218 562 2222
rect 582 2198 586 2202
rect 566 2188 570 2192
rect 550 2168 554 2172
rect 550 2158 554 2162
rect 510 2148 514 2152
rect 558 2148 562 2152
rect 518 2108 522 2112
rect 518 2088 522 2092
rect 526 2068 530 2072
rect 502 2028 506 2032
rect 510 2008 514 2012
rect 526 2008 530 2012
rect 482 2003 486 2007
rect 489 2003 493 2007
rect 502 1998 506 2002
rect 478 1978 482 1982
rect 478 1928 482 1932
rect 470 1918 474 1922
rect 502 1908 506 1912
rect 550 2088 554 2092
rect 678 2308 682 2312
rect 662 2278 666 2282
rect 710 2318 714 2322
rect 790 2378 794 2382
rect 774 2368 778 2372
rect 782 2348 786 2352
rect 798 2348 802 2352
rect 870 2458 874 2462
rect 878 2458 882 2462
rect 838 2438 842 2442
rect 854 2418 858 2422
rect 854 2378 858 2382
rect 822 2358 826 2362
rect 910 2468 914 2472
rect 934 2468 938 2472
rect 902 2458 906 2462
rect 918 2458 922 2462
rect 886 2448 890 2452
rect 926 2448 930 2452
rect 886 2378 890 2382
rect 950 2538 954 2542
rect 998 2538 1002 2542
rect 1038 2538 1042 2542
rect 1070 2538 1074 2542
rect 1094 2540 1098 2544
rect 1126 2538 1130 2542
rect 1150 2538 1154 2542
rect 1174 2538 1178 2542
rect 958 2528 962 2532
rect 1030 2508 1034 2512
rect 994 2503 998 2507
rect 1001 2503 1005 2507
rect 982 2488 986 2492
rect 1110 2518 1114 2522
rect 1062 2498 1066 2502
rect 1126 2528 1130 2532
rect 1238 2598 1242 2602
rect 1406 2838 1410 2842
rect 1390 2808 1394 2812
rect 1398 2758 1402 2762
rect 1358 2728 1362 2732
rect 1334 2708 1338 2712
rect 1350 2708 1354 2712
rect 1286 2588 1290 2592
rect 1318 2648 1322 2652
rect 1318 2608 1322 2612
rect 1310 2598 1314 2602
rect 1334 2588 1338 2592
rect 1310 2578 1314 2582
rect 1302 2568 1306 2572
rect 1398 2728 1402 2732
rect 1462 2878 1466 2882
rect 1514 3003 1518 3007
rect 1521 3003 1525 3007
rect 1550 3298 1554 3302
rect 1598 3298 1602 3302
rect 1646 3298 1650 3302
rect 1670 3298 1674 3302
rect 1638 3288 1642 3292
rect 1670 3288 1674 3292
rect 1590 3278 1594 3282
rect 1574 3268 1578 3272
rect 1638 3268 1642 3272
rect 1654 3268 1658 3272
rect 1566 3258 1570 3262
rect 1542 3238 1546 3242
rect 1638 3248 1642 3252
rect 1574 3238 1578 3242
rect 1598 3218 1602 3222
rect 1566 3178 1570 3182
rect 1726 3298 1730 3302
rect 1702 3278 1706 3282
rect 1702 3258 1706 3262
rect 1734 3258 1738 3262
rect 1686 3248 1690 3252
rect 1678 3198 1682 3202
rect 1678 3188 1682 3192
rect 1598 3168 1602 3172
rect 1670 3148 1674 3152
rect 1670 3138 1674 3142
rect 1542 3098 1546 3102
rect 1582 3088 1586 3092
rect 1590 3078 1594 3082
rect 1550 3048 1554 3052
rect 1566 3038 1570 3042
rect 1550 3018 1554 3022
rect 1566 2998 1570 3002
rect 1558 2988 1562 2992
rect 1494 2958 1498 2962
rect 1502 2958 1506 2962
rect 1518 2958 1522 2962
rect 1534 2958 1538 2962
rect 1582 3048 1586 3052
rect 1582 3018 1586 3022
rect 1574 2938 1578 2942
rect 1510 2918 1514 2922
rect 1478 2868 1482 2872
rect 1478 2858 1482 2862
rect 1502 2858 1506 2862
rect 1430 2838 1434 2842
rect 1526 2848 1530 2852
rect 1514 2803 1518 2807
rect 1521 2803 1525 2807
rect 1526 2788 1530 2792
rect 1462 2758 1466 2762
rect 1430 2748 1434 2752
rect 1454 2748 1458 2752
rect 1422 2738 1426 2742
rect 1414 2708 1418 2712
rect 1406 2688 1410 2692
rect 1382 2678 1386 2682
rect 1422 2668 1426 2672
rect 1414 2648 1418 2652
rect 1374 2638 1378 2642
rect 1350 2578 1354 2582
rect 1358 2558 1362 2562
rect 1318 2548 1322 2552
rect 1366 2548 1370 2552
rect 1318 2538 1322 2542
rect 1366 2538 1370 2542
rect 1222 2528 1226 2532
rect 1198 2518 1202 2522
rect 1174 2508 1178 2512
rect 1126 2498 1130 2502
rect 1054 2488 1058 2492
rect 1118 2488 1122 2492
rect 1062 2478 1066 2482
rect 1006 2468 1010 2472
rect 1038 2468 1042 2472
rect 1166 2488 1170 2492
rect 1158 2468 1162 2472
rect 998 2458 1002 2462
rect 1078 2458 1082 2462
rect 1134 2458 1138 2462
rect 1158 2458 1162 2462
rect 950 2448 954 2452
rect 966 2438 970 2442
rect 974 2438 978 2442
rect 966 2418 970 2422
rect 918 2378 922 2382
rect 910 2368 914 2372
rect 902 2358 906 2362
rect 862 2348 866 2352
rect 766 2338 770 2342
rect 790 2338 794 2342
rect 822 2338 826 2342
rect 830 2338 834 2342
rect 854 2328 858 2332
rect 726 2318 730 2322
rect 734 2318 738 2322
rect 766 2318 770 2322
rect 806 2318 810 2322
rect 694 2308 698 2312
rect 822 2288 826 2292
rect 758 2278 762 2282
rect 798 2278 802 2282
rect 686 2268 690 2272
rect 766 2268 770 2272
rect 710 2258 714 2262
rect 686 2248 690 2252
rect 750 2248 754 2252
rect 662 2238 666 2242
rect 694 2238 698 2242
rect 846 2278 850 2282
rect 870 2318 874 2322
rect 894 2348 898 2352
rect 910 2348 914 2352
rect 942 2358 946 2362
rect 950 2358 954 2362
rect 1054 2448 1058 2452
rect 998 2438 1002 2442
rect 1038 2438 1042 2442
rect 990 2408 994 2412
rect 982 2398 986 2402
rect 1014 2408 1018 2412
rect 1006 2348 1010 2352
rect 1030 2398 1034 2402
rect 1046 2398 1050 2402
rect 974 2338 978 2342
rect 854 2268 858 2272
rect 878 2268 882 2272
rect 782 2228 786 2232
rect 758 2218 762 2222
rect 726 2208 730 2212
rect 654 2198 658 2202
rect 718 2198 722 2202
rect 726 2198 730 2202
rect 638 2168 642 2172
rect 678 2168 682 2172
rect 590 2158 594 2162
rect 598 2148 602 2152
rect 622 2148 626 2152
rect 566 2128 570 2132
rect 566 2118 570 2122
rect 606 2118 610 2122
rect 550 2058 554 2062
rect 574 2108 578 2112
rect 590 2098 594 2102
rect 606 2068 610 2072
rect 630 2128 634 2132
rect 622 2098 626 2102
rect 630 2098 634 2102
rect 798 2198 802 2202
rect 822 2168 826 2172
rect 926 2298 930 2302
rect 918 2268 922 2272
rect 1046 2328 1050 2332
rect 958 2308 962 2312
rect 1014 2308 1018 2312
rect 994 2303 998 2307
rect 1001 2303 1005 2307
rect 934 2288 938 2292
rect 998 2288 1002 2292
rect 950 2278 954 2282
rect 910 2258 914 2262
rect 1006 2238 1010 2242
rect 974 2228 978 2232
rect 886 2198 890 2202
rect 894 2198 898 2202
rect 918 2188 922 2192
rect 854 2168 858 2172
rect 894 2168 898 2172
rect 726 2148 730 2152
rect 750 2148 754 2152
rect 774 2148 778 2152
rect 798 2148 802 2152
rect 838 2148 842 2152
rect 686 2138 690 2142
rect 654 2128 658 2132
rect 702 2128 706 2132
rect 710 2128 714 2132
rect 726 2128 730 2132
rect 758 2128 762 2132
rect 646 2118 650 2122
rect 686 2118 690 2122
rect 638 2078 642 2082
rect 638 2068 642 2072
rect 590 2058 594 2062
rect 614 2058 618 2062
rect 654 2058 658 2062
rect 686 2078 690 2082
rect 678 2068 682 2072
rect 534 1998 538 2002
rect 566 1988 570 1992
rect 534 1978 538 1982
rect 550 1978 554 1982
rect 526 1958 530 1962
rect 558 1968 562 1972
rect 558 1938 562 1942
rect 526 1928 530 1932
rect 534 1928 538 1932
rect 526 1908 530 1912
rect 486 1878 490 1882
rect 422 1818 426 1822
rect 462 1848 466 1852
rect 534 1848 538 1852
rect 518 1838 522 1842
rect 526 1828 530 1832
rect 482 1803 486 1807
rect 489 1803 493 1807
rect 470 1798 474 1802
rect 438 1768 442 1772
rect 454 1768 458 1772
rect 422 1748 426 1752
rect 366 1738 370 1742
rect 430 1738 434 1742
rect 406 1728 410 1732
rect 438 1718 442 1722
rect 382 1708 386 1712
rect 390 1678 394 1682
rect 358 1668 362 1672
rect 366 1668 370 1672
rect 438 1668 442 1672
rect 422 1658 426 1662
rect 334 1648 338 1652
rect 318 1638 322 1642
rect 310 1618 314 1622
rect 294 1598 298 1602
rect 318 1598 322 1602
rect 334 1598 338 1602
rect 286 1568 290 1572
rect 310 1568 314 1572
rect 286 1528 290 1532
rect 294 1528 298 1532
rect 318 1538 322 1542
rect 310 1508 314 1512
rect 302 1468 306 1472
rect 286 1458 290 1462
rect 222 1438 226 1442
rect 230 1438 234 1442
rect 262 1408 266 1412
rect 230 1388 234 1392
rect 238 1368 242 1372
rect 254 1348 258 1352
rect 254 1338 258 1342
rect 198 1278 202 1282
rect 190 1268 194 1272
rect 190 1258 194 1262
rect 198 1258 202 1262
rect 190 1248 194 1252
rect 198 1238 202 1242
rect 246 1328 250 1332
rect 262 1328 266 1332
rect 254 1318 258 1322
rect 214 1268 218 1272
rect 350 1628 354 1632
rect 358 1568 362 1572
rect 342 1518 346 1522
rect 326 1508 330 1512
rect 350 1508 354 1512
rect 342 1478 346 1482
rect 326 1458 330 1462
rect 318 1448 322 1452
rect 358 1458 362 1462
rect 350 1428 354 1432
rect 310 1388 314 1392
rect 302 1368 306 1372
rect 254 1278 258 1282
rect 278 1278 282 1282
rect 342 1378 346 1382
rect 318 1368 322 1372
rect 430 1648 434 1652
rect 454 1738 458 1742
rect 486 1738 490 1742
rect 558 1878 562 1882
rect 598 2038 602 2042
rect 614 2008 618 2012
rect 590 1988 594 1992
rect 622 1988 626 1992
rect 654 2038 658 2042
rect 662 2038 666 2042
rect 654 2008 658 2012
rect 662 1988 666 1992
rect 710 2068 714 2072
rect 750 2108 754 2112
rect 758 2108 762 2112
rect 758 2088 762 2092
rect 766 2088 770 2092
rect 750 2078 754 2082
rect 686 2038 690 2042
rect 694 2028 698 2032
rect 694 1978 698 1982
rect 582 1958 586 1962
rect 646 1958 650 1962
rect 662 1958 666 1962
rect 582 1948 586 1952
rect 606 1948 610 1952
rect 638 1948 642 1952
rect 646 1948 650 1952
rect 718 2038 722 2042
rect 742 2058 746 2062
rect 958 2198 962 2202
rect 942 2168 946 2172
rect 982 2168 986 2172
rect 950 2158 954 2162
rect 806 2138 810 2142
rect 822 2138 826 2142
rect 862 2138 866 2142
rect 886 2138 890 2142
rect 934 2138 938 2142
rect 982 2138 986 2142
rect 806 2128 810 2132
rect 798 2098 802 2102
rect 790 2088 794 2092
rect 774 2048 778 2052
rect 742 2028 746 2032
rect 758 2028 762 2032
rect 734 1988 738 1992
rect 734 1978 738 1982
rect 710 1948 714 1952
rect 630 1938 634 1942
rect 646 1938 650 1942
rect 662 1938 666 1942
rect 574 1908 578 1912
rect 590 1878 594 1882
rect 614 1878 618 1882
rect 582 1868 586 1872
rect 614 1858 618 1862
rect 590 1848 594 1852
rect 550 1828 554 1832
rect 590 1828 594 1832
rect 542 1768 546 1772
rect 526 1748 530 1752
rect 534 1738 538 1742
rect 502 1728 506 1732
rect 510 1728 514 1732
rect 478 1698 482 1702
rect 534 1718 538 1722
rect 454 1658 458 1662
rect 510 1658 514 1662
rect 534 1698 538 1702
rect 566 1788 570 1792
rect 558 1718 562 1722
rect 606 1818 610 1822
rect 598 1798 602 1802
rect 646 1928 650 1932
rect 638 1918 642 1922
rect 630 1908 634 1912
rect 622 1778 626 1782
rect 766 1988 770 1992
rect 790 1988 794 1992
rect 774 1968 778 1972
rect 782 1968 786 1972
rect 838 2098 842 2102
rect 838 2088 842 2092
rect 854 2078 858 2082
rect 918 2118 922 2122
rect 1054 2298 1058 2302
rect 1046 2278 1050 2282
rect 1054 2278 1058 2282
rect 1070 2408 1074 2412
rect 1062 2268 1066 2272
rect 1094 2448 1098 2452
rect 1118 2448 1122 2452
rect 1142 2438 1146 2442
rect 1126 2398 1130 2402
rect 1150 2378 1154 2382
rect 1110 2368 1114 2372
rect 1118 2368 1122 2372
rect 1142 2368 1146 2372
rect 1110 2348 1114 2352
rect 1094 2338 1098 2342
rect 1102 2278 1106 2282
rect 1086 2258 1090 2262
rect 1078 2198 1082 2202
rect 1014 2168 1018 2172
rect 1054 2168 1058 2172
rect 1070 2168 1074 2172
rect 1102 2208 1106 2212
rect 1094 2168 1098 2172
rect 1206 2478 1210 2482
rect 1182 2438 1186 2442
rect 1166 2408 1170 2412
rect 1182 2408 1186 2412
rect 1158 2368 1162 2372
rect 1190 2368 1194 2372
rect 1254 2498 1258 2502
rect 1246 2488 1250 2492
rect 1254 2478 1258 2482
rect 1238 2468 1242 2472
rect 1230 2458 1234 2462
rect 1238 2458 1242 2462
rect 1262 2458 1266 2462
rect 1230 2448 1234 2452
rect 1286 2508 1290 2512
rect 1358 2508 1362 2512
rect 1326 2498 1330 2502
rect 1326 2488 1330 2492
rect 1294 2478 1298 2482
rect 1302 2468 1306 2472
rect 1374 2498 1378 2502
rect 1374 2468 1378 2472
rect 1406 2578 1410 2582
rect 1390 2568 1394 2572
rect 1446 2708 1450 2712
rect 1462 2728 1466 2732
rect 1510 2738 1514 2742
rect 1502 2728 1506 2732
rect 1470 2708 1474 2712
rect 1470 2688 1474 2692
rect 1550 2918 1554 2922
rect 1598 2928 1602 2932
rect 1566 2908 1570 2912
rect 1566 2888 1570 2892
rect 1582 2888 1586 2892
rect 1542 2878 1546 2882
rect 1574 2868 1578 2872
rect 1574 2788 1578 2792
rect 1534 2768 1538 2772
rect 1542 2768 1546 2772
rect 1574 2768 1578 2772
rect 1542 2758 1546 2762
rect 1542 2748 1546 2752
rect 1534 2688 1538 2692
rect 1526 2678 1530 2682
rect 1454 2658 1458 2662
rect 1486 2658 1490 2662
rect 1502 2658 1506 2662
rect 1566 2738 1570 2742
rect 1646 3108 1650 3112
rect 1662 3118 1666 3122
rect 1654 3098 1658 3102
rect 1790 3268 1794 3272
rect 1822 3258 1826 3262
rect 1806 3248 1810 3252
rect 1766 3228 1770 3232
rect 1742 3178 1746 3182
rect 1686 3168 1690 3172
rect 1774 3168 1778 3172
rect 1822 3168 1826 3172
rect 1686 3158 1690 3162
rect 1726 3158 1730 3162
rect 1694 3148 1698 3152
rect 1726 3148 1730 3152
rect 1734 3148 1738 3152
rect 1766 3148 1770 3152
rect 1782 3148 1786 3152
rect 1822 3148 1826 3152
rect 1718 3138 1722 3142
rect 1734 3138 1738 3142
rect 1694 3128 1698 3132
rect 1806 3128 1810 3132
rect 1678 3118 1682 3122
rect 1638 3088 1642 3092
rect 1662 3088 1666 3092
rect 1710 3088 1714 3092
rect 1622 3078 1626 3082
rect 1614 3068 1618 3072
rect 1630 3068 1634 3072
rect 1678 3068 1682 3072
rect 1630 3048 1634 3052
rect 1654 3048 1658 3052
rect 1622 3038 1626 3042
rect 1646 3038 1650 3042
rect 1686 2958 1690 2962
rect 1702 3058 1706 3062
rect 1702 3018 1706 3022
rect 1694 2948 1698 2952
rect 1622 2928 1626 2932
rect 1630 2928 1634 2932
rect 1654 2928 1658 2932
rect 1654 2918 1658 2922
rect 1606 2908 1610 2912
rect 1614 2908 1618 2912
rect 1646 2908 1650 2912
rect 1630 2878 1634 2882
rect 1734 3038 1738 3042
rect 1726 3008 1730 3012
rect 1726 2968 1730 2972
rect 1758 3118 1762 3122
rect 1806 3108 1810 3112
rect 1814 3108 1818 3112
rect 1766 3098 1770 3102
rect 1742 2968 1746 2972
rect 1846 3258 1850 3262
rect 1854 3218 1858 3222
rect 1854 3168 1858 3172
rect 1846 3158 1850 3162
rect 1846 3128 1850 3132
rect 1838 3108 1842 3112
rect 1830 3098 1834 3102
rect 1814 3078 1818 3082
rect 1790 3068 1794 3072
rect 1822 3068 1826 3072
rect 1878 3248 1882 3252
rect 1870 3178 1874 3182
rect 1870 3128 1874 3132
rect 1846 3038 1850 3042
rect 1862 3038 1866 3042
rect 1862 3018 1866 3022
rect 1822 2998 1826 3002
rect 1830 2998 1834 3002
rect 1774 2988 1778 2992
rect 1774 2978 1778 2982
rect 1782 2958 1786 2962
rect 1718 2908 1722 2912
rect 1726 2878 1730 2882
rect 1742 2928 1746 2932
rect 1766 2928 1770 2932
rect 1750 2878 1754 2882
rect 1766 2878 1770 2882
rect 1838 2988 1842 2992
rect 1878 3118 1882 3122
rect 1950 3298 1954 3302
rect 1918 3278 1922 3282
rect 1894 3258 1898 3262
rect 1902 3248 1906 3252
rect 1958 3259 1962 3263
rect 1934 3228 1938 3232
rect 1902 3168 1906 3172
rect 2026 3303 2030 3307
rect 2033 3303 2037 3307
rect 1990 3298 1994 3302
rect 2230 3298 2234 3302
rect 2246 3298 2250 3302
rect 2262 3298 2266 3302
rect 2118 3288 2122 3292
rect 2182 3288 2186 3292
rect 2238 3288 2242 3292
rect 2254 3288 2258 3292
rect 2014 3278 2018 3282
rect 2070 3278 2074 3282
rect 2086 3278 2090 3282
rect 2142 3278 2146 3282
rect 2030 3258 2034 3262
rect 2054 3258 2058 3262
rect 2078 3258 2082 3262
rect 2110 3258 2114 3262
rect 2262 3278 2266 3282
rect 2142 3258 2146 3262
rect 2158 3258 2162 3262
rect 2206 3258 2210 3262
rect 2230 3258 2234 3262
rect 2134 3218 2138 3222
rect 1974 3198 1978 3202
rect 1958 3178 1962 3182
rect 2198 3238 2202 3242
rect 2222 3228 2226 3232
rect 2254 3228 2258 3232
rect 2158 3178 2162 3182
rect 2166 3168 2170 3172
rect 2230 3168 2234 3172
rect 2246 3168 2250 3172
rect 1902 3158 1906 3162
rect 1934 3158 1938 3162
rect 2030 3158 2034 3162
rect 2110 3158 2114 3162
rect 2134 3158 2138 3162
rect 1966 3148 1970 3152
rect 2014 3148 2018 3152
rect 2054 3147 2058 3151
rect 2150 3148 2154 3152
rect 2222 3158 2226 3162
rect 1974 3138 1978 3142
rect 2118 3138 2122 3142
rect 2158 3138 2162 3142
rect 2278 3298 2282 3302
rect 2294 3298 2298 3302
rect 2470 3298 2474 3302
rect 2526 3298 2530 3302
rect 2630 3298 2634 3302
rect 2662 3298 2666 3302
rect 2398 3288 2402 3292
rect 2478 3288 2482 3292
rect 2486 3288 2490 3292
rect 2646 3288 2650 3292
rect 2398 3278 2402 3282
rect 2502 3278 2506 3282
rect 2630 3278 2634 3282
rect 2638 3278 2642 3282
rect 2670 3278 2674 3282
rect 2374 3268 2378 3272
rect 2302 3258 2306 3262
rect 2286 3238 2290 3242
rect 2454 3268 2458 3272
rect 2430 3258 2434 3262
rect 2510 3258 2514 3262
rect 2438 3238 2442 3242
rect 2334 3218 2338 3222
rect 2358 3218 2362 3222
rect 2446 3208 2450 3212
rect 2526 3268 2530 3272
rect 2694 3268 2698 3272
rect 2558 3258 2562 3262
rect 2526 3248 2530 3252
rect 2478 3168 2482 3172
rect 2486 3168 2490 3172
rect 2294 3158 2298 3162
rect 2326 3158 2330 3162
rect 2334 3158 2338 3162
rect 2422 3158 2426 3162
rect 2470 3158 2474 3162
rect 2006 3128 2010 3132
rect 2126 3128 2130 3132
rect 2166 3128 2170 3132
rect 2190 3128 2194 3132
rect 2206 3128 2210 3132
rect 1998 3118 2002 3122
rect 1894 3098 1898 3102
rect 1886 3068 1890 3072
rect 2134 3108 2138 3112
rect 2026 3103 2030 3107
rect 2033 3103 2037 3107
rect 2046 3098 2050 3102
rect 1950 3088 1954 3092
rect 1990 3088 1994 3092
rect 2006 3088 2010 3092
rect 1926 3078 1930 3082
rect 2166 3098 2170 3102
rect 2142 3088 2146 3092
rect 2094 3078 2098 3082
rect 2158 3078 2162 3082
rect 1918 3068 1922 3072
rect 2006 3068 2010 3072
rect 2062 3068 2066 3072
rect 2086 3068 2090 3072
rect 2110 3068 2114 3072
rect 2150 3068 2154 3072
rect 1902 3028 1906 3032
rect 1886 2988 1890 2992
rect 1838 2978 1842 2982
rect 1870 2978 1874 2982
rect 1862 2958 1866 2962
rect 1830 2938 1834 2942
rect 1790 2928 1794 2932
rect 1806 2918 1810 2922
rect 1894 2968 1898 2972
rect 2070 3058 2074 3062
rect 2102 3058 2106 3062
rect 2126 3058 2130 3062
rect 1982 3048 1986 3052
rect 2014 3048 2018 3052
rect 1950 3038 1954 3042
rect 1974 3038 1978 3042
rect 2046 3038 2050 3042
rect 1886 2958 1890 2962
rect 1854 2938 1858 2942
rect 1878 2938 1882 2942
rect 1870 2928 1874 2932
rect 1838 2908 1842 2912
rect 1870 2908 1874 2912
rect 1822 2898 1826 2902
rect 1838 2898 1842 2902
rect 1982 3028 1986 3032
rect 2102 3048 2106 3052
rect 2078 3028 2082 3032
rect 2118 3048 2122 3052
rect 2110 3028 2114 3032
rect 2158 3028 2162 3032
rect 1990 2978 1994 2982
rect 2046 2978 2050 2982
rect 2062 2968 2066 2972
rect 2046 2958 2050 2962
rect 2070 2958 2074 2962
rect 2150 2958 2154 2962
rect 1894 2938 1898 2942
rect 1918 2938 1922 2942
rect 1934 2938 1938 2942
rect 1990 2938 1994 2942
rect 1998 2938 2002 2942
rect 2014 2938 2018 2942
rect 2062 2948 2066 2952
rect 1894 2918 1898 2922
rect 1918 2908 1922 2912
rect 1934 2898 1938 2902
rect 1822 2878 1826 2882
rect 1854 2878 1858 2882
rect 1870 2878 1874 2882
rect 1654 2868 1658 2872
rect 1718 2868 1722 2872
rect 1734 2868 1738 2872
rect 1774 2868 1778 2872
rect 1638 2858 1642 2862
rect 1614 2838 1618 2842
rect 1662 2838 1666 2842
rect 1590 2808 1594 2812
rect 1638 2808 1642 2812
rect 1598 2758 1602 2762
rect 1630 2758 1634 2762
rect 1630 2738 1634 2742
rect 1662 2738 1666 2742
rect 1582 2728 1586 2732
rect 1574 2718 1578 2722
rect 1638 2728 1642 2732
rect 1654 2728 1658 2732
rect 1606 2718 1610 2722
rect 1646 2718 1650 2722
rect 1590 2678 1594 2682
rect 1614 2708 1618 2712
rect 1630 2708 1634 2712
rect 1566 2668 1570 2672
rect 1598 2668 1602 2672
rect 1622 2668 1626 2672
rect 1574 2658 1578 2662
rect 1542 2648 1546 2652
rect 1558 2648 1562 2652
rect 1598 2648 1602 2652
rect 1526 2638 1530 2642
rect 1582 2638 1586 2642
rect 1454 2598 1458 2602
rect 1430 2588 1434 2592
rect 1478 2588 1482 2592
rect 1422 2568 1426 2572
rect 1550 2608 1554 2612
rect 1514 2603 1518 2607
rect 1521 2603 1525 2607
rect 1574 2598 1578 2602
rect 1550 2588 1554 2592
rect 1558 2588 1562 2592
rect 1526 2558 1530 2562
rect 1438 2548 1442 2552
rect 1454 2548 1458 2552
rect 1470 2548 1474 2552
rect 1518 2548 1522 2552
rect 1406 2528 1410 2532
rect 1422 2528 1426 2532
rect 1406 2488 1410 2492
rect 1622 2648 1626 2652
rect 1614 2608 1618 2612
rect 1590 2598 1594 2602
rect 1534 2548 1538 2552
rect 1558 2548 1562 2552
rect 1622 2548 1626 2552
rect 1550 2538 1554 2542
rect 1566 2538 1570 2542
rect 1470 2528 1474 2532
rect 1518 2528 1522 2532
rect 1454 2518 1458 2522
rect 1478 2508 1482 2512
rect 1446 2498 1450 2502
rect 1470 2498 1474 2502
rect 1454 2488 1458 2492
rect 1414 2478 1418 2482
rect 1462 2478 1466 2482
rect 1430 2468 1434 2472
rect 1206 2438 1210 2442
rect 1214 2398 1218 2402
rect 1246 2398 1250 2402
rect 1262 2398 1266 2402
rect 1214 2368 1218 2372
rect 1230 2348 1234 2352
rect 1254 2348 1258 2352
rect 1134 2338 1138 2342
rect 1198 2338 1202 2342
rect 1246 2338 1250 2342
rect 1166 2328 1170 2332
rect 1142 2298 1146 2302
rect 1118 2238 1122 2242
rect 1174 2298 1178 2302
rect 1174 2288 1178 2292
rect 1166 2278 1170 2282
rect 1182 2278 1186 2282
rect 1222 2308 1226 2312
rect 1222 2298 1226 2302
rect 1238 2298 1242 2302
rect 1190 2268 1194 2272
rect 1142 2248 1146 2252
rect 1150 2238 1154 2242
rect 1206 2238 1210 2242
rect 1134 2228 1138 2232
rect 1190 2228 1194 2232
rect 1214 2228 1218 2232
rect 1126 2198 1130 2202
rect 1166 2198 1170 2202
rect 1166 2168 1170 2172
rect 1198 2158 1202 2162
rect 1230 2278 1234 2282
rect 1286 2458 1290 2462
rect 1278 2378 1282 2382
rect 1294 2448 1298 2452
rect 1382 2448 1386 2452
rect 1286 2358 1290 2362
rect 1286 2298 1290 2302
rect 1278 2288 1282 2292
rect 1246 2238 1250 2242
rect 1262 2278 1266 2282
rect 1270 2278 1274 2282
rect 1326 2438 1330 2442
rect 1390 2438 1394 2442
rect 1302 2408 1306 2412
rect 1406 2458 1410 2462
rect 1414 2458 1418 2462
rect 1398 2408 1402 2412
rect 1326 2398 1330 2402
rect 1374 2398 1378 2402
rect 1374 2378 1378 2382
rect 1342 2368 1346 2372
rect 1398 2358 1402 2362
rect 1302 2348 1306 2352
rect 1334 2348 1338 2352
rect 1350 2348 1354 2352
rect 1406 2348 1410 2352
rect 1358 2328 1362 2332
rect 1326 2318 1330 2322
rect 1294 2268 1298 2272
rect 1294 2248 1298 2252
rect 1342 2298 1346 2302
rect 1350 2278 1354 2282
rect 1398 2288 1402 2292
rect 1382 2268 1386 2272
rect 1334 2248 1338 2252
rect 1278 2238 1282 2242
rect 1254 2218 1258 2222
rect 1230 2188 1234 2192
rect 1502 2498 1506 2502
rect 1494 2468 1498 2472
rect 1654 2678 1658 2682
rect 1718 2848 1722 2852
rect 1702 2828 1706 2832
rect 1702 2818 1706 2822
rect 1734 2858 1738 2862
rect 1782 2858 1786 2862
rect 1678 2808 1682 2812
rect 1726 2808 1730 2812
rect 1694 2768 1698 2772
rect 1702 2758 1706 2762
rect 1670 2718 1674 2722
rect 1670 2678 1674 2682
rect 1646 2668 1650 2672
rect 1694 2688 1698 2692
rect 1750 2848 1754 2852
rect 1766 2848 1770 2852
rect 1782 2848 1786 2852
rect 1814 2848 1818 2852
rect 1750 2838 1754 2842
rect 1806 2838 1810 2842
rect 1806 2808 1810 2812
rect 1806 2768 1810 2772
rect 1822 2768 1826 2772
rect 1790 2758 1794 2762
rect 1742 2748 1746 2752
rect 1710 2728 1714 2732
rect 1734 2728 1738 2732
rect 1726 2688 1730 2692
rect 1678 2668 1682 2672
rect 1686 2668 1690 2672
rect 1718 2668 1722 2672
rect 1774 2718 1778 2722
rect 1782 2708 1786 2712
rect 1750 2678 1754 2682
rect 1782 2678 1786 2682
rect 1758 2668 1762 2672
rect 1806 2728 1810 2732
rect 1798 2718 1802 2722
rect 1806 2678 1810 2682
rect 1846 2858 1850 2862
rect 1854 2858 1858 2862
rect 1902 2848 1906 2852
rect 1902 2828 1906 2832
rect 1870 2768 1874 2772
rect 1854 2758 1858 2762
rect 1878 2758 1882 2762
rect 1862 2748 1866 2752
rect 1854 2738 1858 2742
rect 1894 2728 1898 2732
rect 1926 2858 1930 2862
rect 1950 2858 1954 2862
rect 1934 2848 1938 2852
rect 1950 2848 1954 2852
rect 2086 2948 2090 2952
rect 2110 2948 2114 2952
rect 2134 2948 2138 2952
rect 2182 3078 2186 3082
rect 2182 3068 2186 3072
rect 2230 3088 2234 3092
rect 2206 3058 2210 3062
rect 2198 3048 2202 3052
rect 2206 3028 2210 3032
rect 2174 2968 2178 2972
rect 2214 2998 2218 3002
rect 2302 3138 2306 3142
rect 2342 3138 2346 3142
rect 2254 3128 2258 3132
rect 2246 3088 2250 3092
rect 2270 3098 2274 3102
rect 2286 3088 2290 3092
rect 2262 3078 2266 3082
rect 2286 3068 2290 3072
rect 2374 3108 2378 3112
rect 2390 3108 2394 3112
rect 2502 3158 2506 3162
rect 2538 3203 2542 3207
rect 2545 3203 2549 3207
rect 2534 3138 2538 3142
rect 2454 3128 2458 3132
rect 2470 3118 2474 3122
rect 2462 3098 2466 3102
rect 2510 3118 2514 3122
rect 2510 3098 2514 3102
rect 2494 3088 2498 3092
rect 2590 3248 2594 3252
rect 2638 3248 2642 3252
rect 2614 3238 2618 3242
rect 2590 3218 2594 3222
rect 2574 3138 2578 3142
rect 2390 3078 2394 3082
rect 2430 3078 2434 3082
rect 2446 3078 2450 3082
rect 2470 3078 2474 3082
rect 2518 3078 2522 3082
rect 2534 3078 2538 3082
rect 2406 3068 2410 3072
rect 2462 3068 2466 3072
rect 2486 3068 2490 3072
rect 2342 3058 2346 3062
rect 2262 3038 2266 3042
rect 2302 3038 2306 3042
rect 2238 2998 2242 3002
rect 2230 2978 2234 2982
rect 2238 2978 2242 2982
rect 2182 2958 2186 2962
rect 2206 2958 2210 2962
rect 2182 2948 2186 2952
rect 2198 2948 2202 2952
rect 2222 2948 2226 2952
rect 2078 2938 2082 2942
rect 2070 2928 2074 2932
rect 1990 2918 1994 2922
rect 2026 2903 2030 2907
rect 2033 2903 2037 2907
rect 1966 2878 1970 2882
rect 1982 2878 1986 2882
rect 1966 2848 1970 2852
rect 1958 2818 1962 2822
rect 1990 2858 1994 2862
rect 1982 2828 1986 2832
rect 2006 2828 2010 2832
rect 1974 2778 1978 2782
rect 1926 2768 1930 2772
rect 1910 2738 1914 2742
rect 1902 2718 1906 2722
rect 1838 2688 1842 2692
rect 1926 2718 1930 2722
rect 1974 2728 1978 2732
rect 1974 2708 1978 2712
rect 1966 2688 1970 2692
rect 1822 2678 1826 2682
rect 1894 2678 1898 2682
rect 1694 2658 1698 2662
rect 1734 2658 1738 2662
rect 1654 2608 1658 2612
rect 1678 2598 1682 2602
rect 1646 2558 1650 2562
rect 1678 2548 1682 2552
rect 1606 2528 1610 2532
rect 1614 2528 1618 2532
rect 1606 2518 1610 2522
rect 1598 2498 1602 2502
rect 1582 2488 1586 2492
rect 1590 2488 1594 2492
rect 1574 2478 1578 2482
rect 1582 2478 1586 2482
rect 1534 2468 1538 2472
rect 1558 2468 1562 2472
rect 1462 2448 1466 2452
rect 1422 2438 1426 2442
rect 1422 2408 1426 2412
rect 1462 2388 1466 2392
rect 1430 2378 1434 2382
rect 1398 2258 1402 2262
rect 1454 2348 1458 2352
rect 1478 2368 1482 2372
rect 1502 2448 1506 2452
rect 1518 2448 1522 2452
rect 1518 2438 1522 2442
rect 1514 2403 1518 2407
rect 1521 2403 1525 2407
rect 1510 2388 1514 2392
rect 1454 2308 1458 2312
rect 1438 2288 1442 2292
rect 1494 2338 1498 2342
rect 1526 2358 1530 2362
rect 1654 2518 1658 2522
rect 1630 2508 1634 2512
rect 1622 2478 1626 2482
rect 1726 2648 1730 2652
rect 1774 2638 1778 2642
rect 1710 2598 1714 2602
rect 1702 2558 1706 2562
rect 1694 2548 1698 2552
rect 1718 2548 1722 2552
rect 1742 2548 1746 2552
rect 1686 2538 1690 2542
rect 1654 2498 1658 2502
rect 1686 2498 1690 2502
rect 1662 2488 1666 2492
rect 1678 2488 1682 2492
rect 1734 2538 1738 2542
rect 1702 2478 1706 2482
rect 1606 2468 1610 2472
rect 1638 2468 1642 2472
rect 1542 2448 1546 2452
rect 1566 2448 1570 2452
rect 1550 2438 1554 2442
rect 1550 2408 1554 2412
rect 1542 2388 1546 2392
rect 1558 2388 1562 2392
rect 1582 2448 1586 2452
rect 1646 2398 1650 2402
rect 1678 2438 1682 2442
rect 1702 2408 1706 2412
rect 1654 2388 1658 2392
rect 1686 2388 1690 2392
rect 1574 2368 1578 2372
rect 1606 2358 1610 2362
rect 1614 2358 1618 2362
rect 1662 2358 1666 2362
rect 1574 2348 1578 2352
rect 1654 2348 1658 2352
rect 1606 2338 1610 2342
rect 1526 2328 1530 2332
rect 1590 2308 1594 2312
rect 1638 2328 1642 2332
rect 1598 2298 1602 2302
rect 1654 2298 1658 2302
rect 1566 2288 1570 2292
rect 1630 2288 1634 2292
rect 1446 2278 1450 2282
rect 1502 2278 1506 2282
rect 1446 2268 1450 2272
rect 1470 2268 1474 2272
rect 1550 2278 1554 2282
rect 1566 2278 1570 2282
rect 1574 2278 1578 2282
rect 1534 2268 1538 2272
rect 1542 2268 1546 2272
rect 1558 2268 1562 2272
rect 1582 2268 1586 2272
rect 1614 2268 1618 2272
rect 1654 2268 1658 2272
rect 1454 2258 1458 2262
rect 1606 2258 1610 2262
rect 1374 2248 1378 2252
rect 1350 2228 1354 2232
rect 1278 2198 1282 2202
rect 1310 2188 1314 2192
rect 1374 2198 1378 2202
rect 1342 2188 1346 2192
rect 1262 2158 1266 2162
rect 1278 2158 1282 2162
rect 1326 2158 1330 2162
rect 998 2148 1002 2152
rect 1110 2148 1114 2152
rect 1118 2148 1122 2152
rect 1150 2148 1154 2152
rect 1190 2148 1194 2152
rect 1222 2148 1226 2152
rect 1254 2148 1258 2152
rect 1278 2148 1282 2152
rect 1334 2148 1338 2152
rect 1062 2138 1066 2142
rect 1110 2138 1114 2142
rect 870 2108 874 2112
rect 838 2058 842 2062
rect 862 2058 866 2062
rect 910 2098 914 2102
rect 950 2088 954 2092
rect 926 2078 930 2082
rect 894 2068 898 2072
rect 902 2058 906 2062
rect 798 1968 802 1972
rect 758 1948 762 1952
rect 766 1938 770 1942
rect 774 1938 778 1942
rect 694 1928 698 1932
rect 742 1928 746 1932
rect 750 1928 754 1932
rect 678 1898 682 1902
rect 646 1858 650 1862
rect 694 1898 698 1902
rect 718 1868 722 1872
rect 622 1748 626 1752
rect 614 1738 618 1742
rect 590 1718 594 1722
rect 582 1708 586 1712
rect 598 1688 602 1692
rect 534 1668 538 1672
rect 550 1668 554 1672
rect 526 1658 530 1662
rect 446 1618 450 1622
rect 390 1608 394 1612
rect 382 1598 386 1602
rect 482 1603 486 1607
rect 489 1603 493 1607
rect 406 1598 410 1602
rect 398 1568 402 1572
rect 422 1568 426 1572
rect 446 1568 450 1572
rect 470 1568 474 1572
rect 534 1638 538 1642
rect 542 1598 546 1602
rect 526 1568 530 1572
rect 502 1548 506 1552
rect 374 1538 378 1542
rect 414 1538 418 1542
rect 446 1538 450 1542
rect 486 1538 490 1542
rect 374 1518 378 1522
rect 374 1478 378 1482
rect 390 1488 394 1492
rect 422 1528 426 1532
rect 446 1518 450 1522
rect 502 1518 506 1522
rect 454 1488 458 1492
rect 422 1478 426 1482
rect 414 1468 418 1472
rect 462 1468 466 1472
rect 414 1458 418 1462
rect 446 1458 450 1462
rect 390 1448 394 1452
rect 398 1448 402 1452
rect 430 1448 434 1452
rect 374 1378 378 1382
rect 414 1438 418 1442
rect 398 1428 402 1432
rect 398 1398 402 1402
rect 358 1358 362 1362
rect 366 1358 370 1362
rect 390 1358 394 1362
rect 318 1348 322 1352
rect 366 1348 370 1352
rect 310 1338 314 1342
rect 326 1338 330 1342
rect 318 1298 322 1302
rect 342 1288 346 1292
rect 422 1368 426 1372
rect 374 1298 378 1302
rect 334 1278 338 1282
rect 350 1278 354 1282
rect 358 1278 362 1282
rect 294 1268 298 1272
rect 318 1268 322 1272
rect 222 1248 226 1252
rect 246 1248 250 1252
rect 214 1238 218 1242
rect 238 1238 242 1242
rect 206 1168 210 1172
rect 198 1148 202 1152
rect 262 1198 266 1202
rect 238 1178 242 1182
rect 222 1168 226 1172
rect 94 1138 98 1142
rect 142 1138 146 1142
rect 182 1138 186 1142
rect 206 1138 210 1142
rect 70 1128 74 1132
rect 86 1088 90 1092
rect 38 1078 42 1082
rect 78 1078 82 1082
rect 14 1048 18 1052
rect 6 968 10 972
rect 30 1038 34 1042
rect 62 1068 66 1072
rect 110 1128 114 1132
rect 134 1128 138 1132
rect 118 1098 122 1102
rect 78 1048 82 1052
rect 134 1068 138 1072
rect 150 1068 154 1072
rect 174 1108 178 1112
rect 254 1118 258 1122
rect 182 1068 186 1072
rect 190 1068 194 1072
rect 118 1058 122 1062
rect 110 1048 114 1052
rect 142 1058 146 1062
rect 150 1048 154 1052
rect 174 1058 178 1062
rect 94 1038 98 1042
rect 118 1038 122 1042
rect 86 1008 90 1012
rect 38 968 42 972
rect 86 968 90 972
rect 78 948 82 952
rect 126 1028 130 1032
rect 126 1018 130 1022
rect 134 1008 138 1012
rect 102 968 106 972
rect 110 948 114 952
rect 30 938 34 942
rect 70 938 74 942
rect 46 908 50 912
rect 14 878 18 882
rect 30 878 34 882
rect 62 878 66 882
rect 14 868 18 872
rect 174 1038 178 1042
rect 158 968 162 972
rect 238 1058 242 1062
rect 190 1018 194 1022
rect 286 1248 290 1252
rect 350 1268 354 1272
rect 318 1238 322 1242
rect 334 1238 338 1242
rect 310 1208 314 1212
rect 318 1208 322 1212
rect 270 1178 274 1182
rect 286 1168 290 1172
rect 318 1178 322 1182
rect 270 1148 274 1152
rect 318 1148 322 1152
rect 390 1298 394 1302
rect 366 1268 370 1272
rect 382 1268 386 1272
rect 374 1248 378 1252
rect 342 1148 346 1152
rect 270 1118 274 1122
rect 206 1038 210 1042
rect 238 968 242 972
rect 294 1068 298 1072
rect 294 1058 298 1062
rect 278 1038 282 1042
rect 342 1078 346 1082
rect 350 1068 354 1072
rect 334 1058 338 1062
rect 350 1058 354 1062
rect 398 1278 402 1282
rect 422 1278 426 1282
rect 398 1268 402 1272
rect 414 1268 418 1272
rect 398 1248 402 1252
rect 398 1188 402 1192
rect 494 1468 498 1472
rect 478 1438 482 1442
rect 454 1428 458 1432
rect 482 1403 486 1407
rect 489 1403 493 1407
rect 494 1388 498 1392
rect 486 1378 490 1382
rect 446 1368 450 1372
rect 438 1358 442 1362
rect 462 1358 466 1362
rect 462 1348 466 1352
rect 454 1338 458 1342
rect 438 1328 442 1332
rect 446 1318 450 1322
rect 454 1288 458 1292
rect 486 1288 490 1292
rect 438 1278 442 1282
rect 446 1268 450 1272
rect 494 1268 498 1272
rect 574 1678 578 1682
rect 558 1598 562 1602
rect 550 1548 554 1552
rect 534 1538 538 1542
rect 582 1668 586 1672
rect 598 1668 602 1672
rect 638 1738 642 1742
rect 662 1758 666 1762
rect 694 1848 698 1852
rect 742 1908 746 1912
rect 774 1908 778 1912
rect 798 1878 802 1882
rect 750 1868 754 1872
rect 766 1868 770 1872
rect 822 1938 826 1942
rect 846 2038 850 2042
rect 854 1948 858 1952
rect 918 2048 922 2052
rect 942 2048 946 2052
rect 886 2038 890 2042
rect 910 1978 914 1982
rect 926 1968 930 1972
rect 994 2103 998 2107
rect 1001 2103 1005 2107
rect 998 2068 1002 2072
rect 982 2058 986 2062
rect 1038 2088 1042 2092
rect 1030 2078 1034 2082
rect 1094 2128 1098 2132
rect 1086 2118 1090 2122
rect 1110 2118 1114 2122
rect 1070 2108 1074 2112
rect 1070 2088 1074 2092
rect 1054 2078 1058 2082
rect 1046 2068 1050 2072
rect 1054 2058 1058 2062
rect 1062 2038 1066 2042
rect 1006 2028 1010 2032
rect 1014 2028 1018 2032
rect 950 1988 954 1992
rect 1046 1988 1050 1992
rect 958 1978 962 1982
rect 1022 1978 1026 1982
rect 966 1968 970 1972
rect 1038 1968 1042 1972
rect 1030 1958 1034 1962
rect 918 1948 922 1952
rect 942 1948 946 1952
rect 966 1948 970 1952
rect 1014 1948 1018 1952
rect 910 1938 914 1942
rect 862 1908 866 1912
rect 886 1928 890 1932
rect 878 1908 882 1912
rect 870 1898 874 1902
rect 822 1878 826 1882
rect 830 1868 834 1872
rect 862 1868 866 1872
rect 758 1858 762 1862
rect 766 1858 770 1862
rect 774 1858 778 1862
rect 814 1858 818 1862
rect 838 1858 842 1862
rect 734 1848 738 1852
rect 678 1748 682 1752
rect 646 1718 650 1722
rect 654 1708 658 1712
rect 678 1708 682 1712
rect 646 1688 650 1692
rect 630 1678 634 1682
rect 710 1768 714 1772
rect 718 1768 722 1772
rect 758 1798 762 1802
rect 702 1748 706 1752
rect 734 1748 738 1752
rect 694 1738 698 1742
rect 718 1738 722 1742
rect 694 1718 698 1722
rect 686 1678 690 1682
rect 638 1668 642 1672
rect 662 1668 666 1672
rect 614 1658 618 1662
rect 630 1658 634 1662
rect 606 1598 610 1602
rect 630 1598 634 1602
rect 598 1588 602 1592
rect 566 1568 570 1572
rect 574 1548 578 1552
rect 590 1548 594 1552
rect 598 1548 602 1552
rect 678 1598 682 1602
rect 670 1578 674 1582
rect 630 1548 634 1552
rect 654 1548 658 1552
rect 574 1528 578 1532
rect 606 1528 610 1532
rect 582 1498 586 1502
rect 598 1478 602 1482
rect 622 1538 626 1542
rect 654 1538 658 1542
rect 558 1468 562 1472
rect 598 1468 602 1472
rect 614 1468 618 1472
rect 518 1458 522 1462
rect 534 1458 538 1462
rect 558 1458 562 1462
rect 598 1458 602 1462
rect 638 1508 642 1512
rect 638 1498 642 1502
rect 550 1448 554 1452
rect 646 1468 650 1472
rect 662 1458 666 1462
rect 598 1448 602 1452
rect 638 1448 642 1452
rect 590 1438 594 1442
rect 622 1438 626 1442
rect 646 1438 650 1442
rect 510 1418 514 1422
rect 526 1368 530 1372
rect 582 1408 586 1412
rect 638 1388 642 1392
rect 606 1378 610 1382
rect 534 1358 538 1362
rect 558 1358 562 1362
rect 566 1358 570 1362
rect 606 1358 610 1362
rect 430 1258 434 1262
rect 422 1248 426 1252
rect 486 1248 490 1252
rect 454 1238 458 1242
rect 446 1188 450 1192
rect 414 1148 418 1152
rect 438 1148 442 1152
rect 398 1138 402 1142
rect 422 1138 426 1142
rect 438 1118 442 1122
rect 470 1208 474 1212
rect 482 1203 486 1207
rect 489 1203 493 1207
rect 502 1198 506 1202
rect 534 1338 538 1342
rect 558 1338 562 1342
rect 582 1338 586 1342
rect 622 1338 626 1342
rect 550 1308 554 1312
rect 598 1328 602 1332
rect 566 1268 570 1272
rect 558 1258 562 1262
rect 518 1218 522 1222
rect 510 1158 514 1162
rect 654 1378 658 1382
rect 646 1318 650 1322
rect 598 1268 602 1272
rect 606 1268 610 1272
rect 622 1268 626 1272
rect 630 1268 634 1272
rect 742 1708 746 1712
rect 710 1678 714 1682
rect 742 1658 746 1662
rect 790 1848 794 1852
rect 806 1808 810 1812
rect 798 1798 802 1802
rect 774 1788 778 1792
rect 798 1788 802 1792
rect 814 1788 818 1792
rect 822 1768 826 1772
rect 774 1748 778 1752
rect 766 1738 770 1742
rect 790 1728 794 1732
rect 798 1698 802 1702
rect 814 1708 818 1712
rect 806 1678 810 1682
rect 782 1658 786 1662
rect 798 1658 802 1662
rect 806 1658 810 1662
rect 750 1648 754 1652
rect 718 1638 722 1642
rect 734 1628 738 1632
rect 758 1628 762 1632
rect 790 1618 794 1622
rect 694 1598 698 1602
rect 726 1578 730 1582
rect 774 1568 778 1572
rect 726 1558 730 1562
rect 846 1728 850 1732
rect 854 1698 858 1702
rect 822 1688 826 1692
rect 846 1668 850 1672
rect 830 1658 834 1662
rect 830 1648 834 1652
rect 942 1928 946 1932
rect 934 1898 938 1902
rect 886 1868 890 1872
rect 918 1868 922 1872
rect 934 1868 938 1872
rect 910 1818 914 1822
rect 934 1828 938 1832
rect 926 1798 930 1802
rect 918 1778 922 1782
rect 918 1768 922 1772
rect 1102 2088 1106 2092
rect 1142 2088 1146 2092
rect 1118 2078 1122 2082
rect 1174 2078 1178 2082
rect 1110 2048 1114 2052
rect 1078 2038 1082 2042
rect 1078 2028 1082 2032
rect 1094 1998 1098 2002
rect 1102 1978 1106 1982
rect 1126 1968 1130 1972
rect 1086 1958 1090 1962
rect 1070 1948 1074 1952
rect 974 1938 978 1942
rect 1102 1938 1106 1942
rect 974 1928 978 1932
rect 994 1903 998 1907
rect 1001 1903 1005 1907
rect 974 1898 978 1902
rect 982 1878 986 1882
rect 990 1868 994 1872
rect 966 1848 970 1852
rect 950 1818 954 1822
rect 958 1808 962 1812
rect 966 1778 970 1782
rect 1030 1848 1034 1852
rect 1014 1788 1018 1792
rect 990 1768 994 1772
rect 1030 1768 1034 1772
rect 1110 1888 1114 1892
rect 1054 1878 1058 1882
rect 1086 1878 1090 1882
rect 1086 1868 1090 1872
rect 1054 1778 1058 1782
rect 1014 1758 1018 1762
rect 1038 1758 1042 1762
rect 870 1738 874 1742
rect 886 1738 890 1742
rect 966 1738 970 1742
rect 1030 1738 1034 1742
rect 918 1728 922 1732
rect 934 1728 938 1732
rect 942 1728 946 1732
rect 958 1728 962 1732
rect 878 1718 882 1722
rect 886 1708 890 1712
rect 910 1708 914 1712
rect 910 1698 914 1702
rect 902 1688 906 1692
rect 870 1668 874 1672
rect 862 1648 866 1652
rect 846 1638 850 1642
rect 814 1608 818 1612
rect 830 1608 834 1612
rect 846 1608 850 1612
rect 798 1578 802 1582
rect 806 1558 810 1562
rect 838 1568 842 1572
rect 694 1538 698 1542
rect 710 1538 714 1542
rect 718 1538 722 1542
rect 686 1518 690 1522
rect 710 1518 714 1522
rect 694 1508 698 1512
rect 702 1478 706 1482
rect 710 1468 714 1472
rect 686 1358 690 1362
rect 694 1358 698 1362
rect 702 1348 706 1352
rect 662 1318 666 1322
rect 662 1298 666 1302
rect 590 1258 594 1262
rect 614 1258 618 1262
rect 638 1258 642 1262
rect 646 1258 650 1262
rect 614 1228 618 1232
rect 646 1228 650 1232
rect 566 1218 570 1222
rect 582 1208 586 1212
rect 550 1188 554 1192
rect 558 1158 562 1162
rect 630 1188 634 1192
rect 534 1148 538 1152
rect 606 1148 610 1152
rect 462 1128 466 1132
rect 454 1108 458 1112
rect 502 1108 506 1112
rect 374 1098 378 1102
rect 430 1098 434 1102
rect 526 1138 530 1142
rect 518 1098 522 1102
rect 534 1098 538 1102
rect 406 1088 410 1092
rect 478 1088 482 1092
rect 462 1078 466 1082
rect 366 1068 370 1072
rect 406 1068 410 1072
rect 470 1068 474 1072
rect 390 1058 394 1062
rect 422 1058 426 1062
rect 438 1058 442 1062
rect 454 1058 458 1062
rect 470 1058 474 1062
rect 350 1038 354 1042
rect 374 1028 378 1032
rect 326 1008 330 1012
rect 302 978 306 982
rect 286 968 290 972
rect 310 968 314 972
rect 182 948 186 952
rect 190 938 194 942
rect 78 868 82 872
rect 110 868 114 872
rect 78 858 82 862
rect 94 858 98 862
rect 54 848 58 852
rect 62 848 66 852
rect 70 838 74 842
rect 54 828 58 832
rect 46 808 50 812
rect 166 928 170 932
rect 182 928 186 932
rect 174 918 178 922
rect 142 908 146 912
rect 134 858 138 862
rect 110 848 114 852
rect 126 848 130 852
rect 166 858 170 862
rect 86 838 90 842
rect 78 748 82 752
rect 46 738 50 742
rect 62 738 66 742
rect 46 728 50 732
rect 54 728 58 732
rect 70 728 74 732
rect 30 708 34 712
rect 22 698 26 702
rect 14 678 18 682
rect 14 658 18 662
rect 38 678 42 682
rect 38 668 42 672
rect 14 548 18 552
rect 70 678 74 682
rect 126 838 130 842
rect 358 978 362 982
rect 222 948 226 952
rect 246 948 250 952
rect 278 948 282 952
rect 286 948 290 952
rect 334 948 338 952
rect 206 928 210 932
rect 214 898 218 902
rect 358 938 362 942
rect 366 938 370 942
rect 254 928 258 932
rect 270 928 274 932
rect 294 918 298 922
rect 310 918 314 922
rect 294 898 298 902
rect 286 888 290 892
rect 254 878 258 882
rect 206 868 210 872
rect 222 868 226 872
rect 198 858 202 862
rect 214 858 218 862
rect 230 858 234 862
rect 182 848 186 852
rect 174 828 178 832
rect 126 808 130 812
rect 150 798 154 802
rect 190 838 194 842
rect 182 788 186 792
rect 350 888 354 892
rect 382 988 386 992
rect 390 948 394 952
rect 398 928 402 932
rect 326 878 330 882
rect 366 878 370 882
rect 318 868 322 872
rect 310 858 314 862
rect 262 838 266 842
rect 238 818 242 822
rect 342 858 346 862
rect 334 818 338 822
rect 350 818 354 822
rect 270 798 274 802
rect 334 778 338 782
rect 206 768 210 772
rect 246 768 250 772
rect 262 768 266 772
rect 318 768 322 772
rect 230 758 234 762
rect 94 738 98 742
rect 110 738 114 742
rect 86 728 90 732
rect 118 718 122 722
rect 110 678 114 682
rect 78 668 82 672
rect 62 648 66 652
rect 94 658 98 662
rect 118 668 122 672
rect 142 718 146 722
rect 446 1038 450 1042
rect 510 1058 514 1062
rect 510 1038 514 1042
rect 526 1038 530 1042
rect 482 1003 486 1007
rect 489 1003 493 1007
rect 526 1008 530 1012
rect 454 988 458 992
rect 438 968 442 972
rect 422 938 426 942
rect 422 908 426 912
rect 398 878 402 882
rect 406 878 410 882
rect 430 898 434 902
rect 566 1118 570 1122
rect 558 1088 562 1092
rect 590 1098 594 1102
rect 590 1068 594 1072
rect 622 1078 626 1082
rect 622 1068 626 1072
rect 550 1058 554 1062
rect 582 1058 586 1062
rect 606 1058 610 1062
rect 582 1038 586 1042
rect 590 1038 594 1042
rect 574 958 578 962
rect 534 948 538 952
rect 550 948 554 952
rect 526 938 530 942
rect 486 928 490 932
rect 478 898 482 902
rect 478 888 482 892
rect 454 878 458 882
rect 486 878 490 882
rect 542 938 546 942
rect 550 938 554 942
rect 606 948 610 952
rect 718 1438 722 1442
rect 750 1538 754 1542
rect 758 1508 762 1512
rect 822 1538 826 1542
rect 750 1478 754 1482
rect 734 1468 738 1472
rect 766 1468 770 1472
rect 758 1448 762 1452
rect 798 1448 802 1452
rect 742 1438 746 1442
rect 774 1438 778 1442
rect 782 1438 786 1442
rect 822 1498 826 1502
rect 822 1488 826 1492
rect 838 1498 842 1502
rect 886 1638 890 1642
rect 862 1568 866 1572
rect 878 1568 882 1572
rect 886 1568 890 1572
rect 894 1568 898 1572
rect 870 1548 874 1552
rect 870 1528 874 1532
rect 854 1508 858 1512
rect 878 1508 882 1512
rect 894 1478 898 1482
rect 870 1468 874 1472
rect 830 1458 834 1462
rect 958 1718 962 1722
rect 926 1708 930 1712
rect 934 1688 938 1692
rect 1054 1728 1058 1732
rect 966 1708 970 1712
rect 926 1668 930 1672
rect 966 1668 970 1672
rect 942 1648 946 1652
rect 918 1578 922 1582
rect 910 1568 914 1572
rect 934 1568 938 1572
rect 918 1548 922 1552
rect 934 1548 938 1552
rect 950 1548 954 1552
rect 934 1528 938 1532
rect 958 1528 962 1532
rect 958 1518 962 1522
rect 918 1508 922 1512
rect 926 1508 930 1512
rect 994 1703 998 1707
rect 1001 1703 1005 1707
rect 1030 1698 1034 1702
rect 1014 1688 1018 1692
rect 1054 1678 1058 1682
rect 1038 1668 1042 1672
rect 1086 1778 1090 1782
rect 1078 1758 1082 1762
rect 1094 1768 1098 1772
rect 1246 2118 1250 2122
rect 1302 2128 1306 2132
rect 1326 2128 1330 2132
rect 1318 2118 1322 2122
rect 1278 2108 1282 2112
rect 1302 2108 1306 2112
rect 1230 2098 1234 2102
rect 1262 2098 1266 2102
rect 1206 2088 1210 2092
rect 1214 2088 1218 2092
rect 1222 2088 1226 2092
rect 1142 2048 1146 2052
rect 1166 2048 1170 2052
rect 1198 2038 1202 2042
rect 1174 1978 1178 1982
rect 1190 1978 1194 1982
rect 1166 1948 1170 1952
rect 1174 1948 1178 1952
rect 1142 1938 1146 1942
rect 1190 1938 1194 1942
rect 1206 1928 1210 1932
rect 1286 2088 1290 2092
rect 1326 2088 1330 2092
rect 1334 2088 1338 2092
rect 1382 2178 1386 2182
rect 1358 2158 1362 2162
rect 1414 2248 1418 2252
rect 1438 2248 1442 2252
rect 1438 2238 1442 2242
rect 1406 2158 1410 2162
rect 1398 2148 1402 2152
rect 1262 2068 1266 2072
rect 1278 2068 1282 2072
rect 1302 2068 1306 2072
rect 1318 2068 1322 2072
rect 1326 2068 1330 2072
rect 1246 2048 1250 2052
rect 1262 1998 1266 2002
rect 1222 1988 1226 1992
rect 1270 1988 1274 1992
rect 1286 1988 1290 1992
rect 1270 1978 1274 1982
rect 1238 1968 1242 1972
rect 1358 2088 1362 2092
rect 1366 2088 1370 2092
rect 1382 2088 1386 2092
rect 1390 2088 1394 2092
rect 1398 2078 1402 2082
rect 1398 2048 1402 2052
rect 1446 2158 1450 2162
rect 1470 2248 1474 2252
rect 1598 2248 1602 2252
rect 1558 2238 1562 2242
rect 1502 2228 1506 2232
rect 1486 2198 1490 2202
rect 1514 2203 1518 2207
rect 1521 2203 1525 2207
rect 1510 2178 1514 2182
rect 1534 2178 1538 2182
rect 1558 2178 1562 2182
rect 1502 2128 1506 2132
rect 1438 2098 1442 2102
rect 1430 2088 1434 2092
rect 1454 2088 1458 2092
rect 1422 2068 1426 2072
rect 1486 2088 1490 2092
rect 1510 2118 1514 2122
rect 1414 2048 1418 2052
rect 1614 2178 1618 2182
rect 1702 2348 1706 2352
rect 1734 2518 1738 2522
rect 1718 2508 1722 2512
rect 1886 2668 1890 2672
rect 1910 2678 1914 2682
rect 1918 2668 1922 2672
rect 1942 2668 1946 2672
rect 1958 2668 1962 2672
rect 1870 2658 1874 2662
rect 1854 2648 1858 2652
rect 1886 2648 1890 2652
rect 1902 2648 1906 2652
rect 1838 2618 1842 2622
rect 1846 2608 1850 2612
rect 1846 2598 1850 2602
rect 1822 2588 1826 2592
rect 1790 2578 1794 2582
rect 1822 2578 1826 2582
rect 1766 2558 1770 2562
rect 1758 2548 1762 2552
rect 1886 2558 1890 2562
rect 1894 2558 1898 2562
rect 1830 2548 1834 2552
rect 1854 2548 1858 2552
rect 1926 2548 1930 2552
rect 1958 2548 1962 2552
rect 1790 2538 1794 2542
rect 1838 2538 1842 2542
rect 1862 2538 1866 2542
rect 1886 2538 1890 2542
rect 1910 2538 1914 2542
rect 1934 2538 1938 2542
rect 1750 2488 1754 2492
rect 1782 2508 1786 2512
rect 1774 2488 1778 2492
rect 1790 2498 1794 2502
rect 1822 2488 1826 2492
rect 1854 2518 1858 2522
rect 1926 2518 1930 2522
rect 1926 2508 1930 2512
rect 1830 2478 1834 2482
rect 1718 2448 1722 2452
rect 1742 2448 1746 2452
rect 1766 2448 1770 2452
rect 1798 2448 1802 2452
rect 1774 2438 1778 2442
rect 1822 2468 1826 2472
rect 1822 2448 1826 2452
rect 1750 2418 1754 2422
rect 1806 2418 1810 2422
rect 1838 2418 1842 2422
rect 1878 2468 1882 2472
rect 1862 2418 1866 2422
rect 1886 2418 1890 2422
rect 1910 2468 1914 2472
rect 1942 2518 1946 2522
rect 1942 2498 1946 2502
rect 1998 2768 2002 2772
rect 1990 2718 1994 2722
rect 2006 2718 2010 2722
rect 2006 2688 2010 2692
rect 1998 2608 2002 2612
rect 1966 2538 1970 2542
rect 1982 2528 1986 2532
rect 1990 2498 1994 2502
rect 2022 2808 2026 2812
rect 2094 2918 2098 2922
rect 2126 2918 2130 2922
rect 2102 2898 2106 2902
rect 2118 2878 2122 2882
rect 2062 2858 2066 2862
rect 2054 2848 2058 2852
rect 2118 2848 2122 2852
rect 2094 2828 2098 2832
rect 2038 2778 2042 2782
rect 2118 2768 2122 2772
rect 2046 2758 2050 2762
rect 2054 2758 2058 2762
rect 2086 2758 2090 2762
rect 2038 2738 2042 2742
rect 2026 2703 2030 2707
rect 2033 2703 2037 2707
rect 2054 2748 2058 2752
rect 2062 2748 2066 2752
rect 2118 2748 2122 2752
rect 2078 2738 2082 2742
rect 2110 2738 2114 2742
rect 2078 2728 2082 2732
rect 2110 2728 2114 2732
rect 2150 2908 2154 2912
rect 2150 2888 2154 2892
rect 2166 2868 2170 2872
rect 2142 2828 2146 2832
rect 2158 2828 2162 2832
rect 2214 2938 2218 2942
rect 2222 2938 2226 2942
rect 2206 2878 2210 2882
rect 2214 2878 2218 2882
rect 2230 2898 2234 2902
rect 2198 2868 2202 2872
rect 2222 2858 2226 2862
rect 2278 2958 2282 2962
rect 2334 2958 2338 2962
rect 2270 2948 2274 2952
rect 2326 2948 2330 2952
rect 2270 2938 2274 2942
rect 2278 2938 2282 2942
rect 2310 2938 2314 2942
rect 2422 3058 2426 3062
rect 2494 3058 2498 3062
rect 2454 3048 2458 3052
rect 2486 3048 2490 3052
rect 2502 3048 2506 3052
rect 2430 3038 2434 3042
rect 2446 3038 2450 3042
rect 2438 3008 2442 3012
rect 2430 2998 2434 3002
rect 2438 2978 2442 2982
rect 2366 2938 2370 2942
rect 2438 2928 2442 2932
rect 2374 2918 2378 2922
rect 2286 2898 2290 2902
rect 2238 2888 2242 2892
rect 2254 2888 2258 2892
rect 2246 2868 2250 2872
rect 2238 2858 2242 2862
rect 2206 2848 2210 2852
rect 2198 2838 2202 2842
rect 2190 2828 2194 2832
rect 2174 2798 2178 2802
rect 2166 2768 2170 2772
rect 2190 2768 2194 2772
rect 2182 2748 2186 2752
rect 2222 2798 2226 2802
rect 2246 2798 2250 2802
rect 2246 2778 2250 2782
rect 2214 2748 2218 2752
rect 2230 2748 2234 2752
rect 2302 2888 2306 2892
rect 2286 2868 2290 2872
rect 2270 2858 2274 2862
rect 2294 2858 2298 2862
rect 2270 2848 2274 2852
rect 2302 2818 2306 2822
rect 2270 2778 2274 2782
rect 2254 2768 2258 2772
rect 2262 2768 2266 2772
rect 2190 2738 2194 2742
rect 2222 2738 2226 2742
rect 2262 2758 2266 2762
rect 2278 2758 2282 2762
rect 2278 2738 2282 2742
rect 2182 2728 2186 2732
rect 2198 2728 2202 2732
rect 2126 2718 2130 2722
rect 2238 2708 2242 2712
rect 2222 2698 2226 2702
rect 2254 2688 2258 2692
rect 2062 2678 2066 2682
rect 2158 2678 2162 2682
rect 2166 2678 2170 2682
rect 2206 2678 2210 2682
rect 2238 2678 2242 2682
rect 2294 2748 2298 2752
rect 2302 2688 2306 2692
rect 2102 2668 2106 2672
rect 2118 2668 2122 2672
rect 2022 2648 2026 2652
rect 2190 2668 2194 2672
rect 2222 2668 2226 2672
rect 2094 2658 2098 2662
rect 2102 2658 2106 2662
rect 2126 2658 2130 2662
rect 2134 2658 2138 2662
rect 2150 2658 2154 2662
rect 2182 2658 2186 2662
rect 2014 2638 2018 2642
rect 2062 2638 2066 2642
rect 2006 2598 2010 2602
rect 2054 2578 2058 2582
rect 2102 2578 2106 2582
rect 2014 2568 2018 2572
rect 2006 2548 2010 2552
rect 2030 2548 2034 2552
rect 2046 2538 2050 2542
rect 2014 2528 2018 2532
rect 2022 2528 2026 2532
rect 2026 2503 2030 2507
rect 2033 2503 2037 2507
rect 1966 2488 1970 2492
rect 1990 2488 1994 2492
rect 2126 2548 2130 2552
rect 2070 2528 2074 2532
rect 2086 2528 2090 2532
rect 2054 2518 2058 2522
rect 2078 2508 2082 2512
rect 2054 2498 2058 2502
rect 2070 2498 2074 2502
rect 1934 2478 1938 2482
rect 1950 2468 1954 2472
rect 1974 2468 1978 2472
rect 1990 2468 1994 2472
rect 2022 2468 2026 2472
rect 2070 2488 2074 2492
rect 2078 2488 2082 2492
rect 2102 2488 2106 2492
rect 2086 2478 2090 2482
rect 2102 2478 2106 2482
rect 2222 2638 2226 2642
rect 2318 2898 2322 2902
rect 2518 3048 2522 3052
rect 2510 3038 2514 3042
rect 2582 3108 2586 3112
rect 2662 3258 2666 3262
rect 2702 3258 2706 3262
rect 2654 3238 2658 3242
rect 2814 3298 2818 3302
rect 2926 3298 2930 3302
rect 2934 3298 2938 3302
rect 2798 3288 2802 3292
rect 2814 3278 2818 3282
rect 2774 3268 2778 3272
rect 2726 3238 2730 3242
rect 2798 3258 2802 3262
rect 2822 3258 2826 3262
rect 2838 3258 2842 3262
rect 2854 3258 2858 3262
rect 2782 3228 2786 3232
rect 2670 3178 2674 3182
rect 2702 3168 2706 3172
rect 2710 3168 2714 3172
rect 2646 3158 2650 3162
rect 2678 3158 2682 3162
rect 2854 3248 2858 3252
rect 2886 3248 2890 3252
rect 2830 3238 2834 3242
rect 2822 3218 2826 3222
rect 2894 3228 2898 3232
rect 2958 3298 2962 3302
rect 3042 3303 3046 3307
rect 3049 3303 3053 3307
rect 3086 3298 3090 3302
rect 2950 3278 2954 3282
rect 2982 3278 2986 3282
rect 2942 3258 2946 3262
rect 2926 3168 2930 3172
rect 2734 3138 2738 3142
rect 2886 3148 2890 3152
rect 2782 3138 2786 3142
rect 2654 3128 2658 3132
rect 2686 3128 2690 3132
rect 2790 3128 2794 3132
rect 2798 3128 2802 3132
rect 2806 3128 2810 3132
rect 2558 3068 2562 3072
rect 2582 3068 2586 3072
rect 2654 3068 2658 3072
rect 2518 3028 2522 3032
rect 2526 3028 2530 3032
rect 2538 3003 2542 3007
rect 2545 3003 2549 3007
rect 2622 3058 2626 3062
rect 2574 3018 2578 3022
rect 2462 2968 2466 2972
rect 2518 2958 2522 2962
rect 2558 2958 2562 2962
rect 2494 2948 2498 2952
rect 2542 2948 2546 2952
rect 2582 2948 2586 2952
rect 2462 2928 2466 2932
rect 2478 2918 2482 2922
rect 2446 2908 2450 2912
rect 2390 2888 2394 2892
rect 2398 2888 2402 2892
rect 2510 2938 2514 2942
rect 2494 2928 2498 2932
rect 2606 2928 2610 2932
rect 2502 2898 2506 2902
rect 2630 3048 2634 3052
rect 2702 3118 2706 3122
rect 2686 3108 2690 3112
rect 2750 3108 2754 3112
rect 2838 3118 2842 3122
rect 2862 3118 2866 3122
rect 2870 3118 2874 3122
rect 2702 3078 2706 3082
rect 2862 3078 2866 3082
rect 2782 3068 2786 3072
rect 2718 3048 2722 3052
rect 2670 3038 2674 3042
rect 2718 3038 2722 3042
rect 2710 2998 2714 3002
rect 2806 3058 2810 3062
rect 2822 3048 2826 3052
rect 3006 3248 3010 3252
rect 3054 3248 3058 3252
rect 3030 3238 3034 3242
rect 2966 3178 2970 3182
rect 3086 3248 3090 3252
rect 3094 3248 3098 3252
rect 3070 3238 3074 3242
rect 3078 3238 3082 3242
rect 2958 3158 2962 3162
rect 2974 3158 2978 3162
rect 3014 3158 3018 3162
rect 2918 3118 2922 3122
rect 2846 3058 2850 3062
rect 2918 3058 2922 3062
rect 2950 3058 2954 3062
rect 2758 3018 2762 3022
rect 2830 3018 2834 3022
rect 2734 2978 2738 2982
rect 2662 2948 2666 2952
rect 2734 2938 2738 2942
rect 2670 2928 2674 2932
rect 2694 2928 2698 2932
rect 2726 2918 2730 2922
rect 2646 2898 2650 2902
rect 2462 2888 2466 2892
rect 2486 2888 2490 2892
rect 2502 2888 2506 2892
rect 2534 2888 2538 2892
rect 2630 2888 2634 2892
rect 2430 2878 2434 2882
rect 2374 2868 2378 2872
rect 2414 2868 2418 2872
rect 2422 2868 2426 2872
rect 2446 2868 2450 2872
rect 2334 2858 2338 2862
rect 2358 2858 2362 2862
rect 2326 2848 2330 2852
rect 2326 2828 2330 2832
rect 2366 2848 2370 2852
rect 2590 2878 2594 2882
rect 2638 2878 2642 2882
rect 2782 2998 2786 3002
rect 2806 3008 2810 3012
rect 2934 2968 2938 2972
rect 2838 2958 2842 2962
rect 2870 2948 2874 2952
rect 2878 2948 2882 2952
rect 2894 2948 2898 2952
rect 2918 2948 2922 2952
rect 2942 2948 2946 2952
rect 2798 2928 2802 2932
rect 2774 2908 2778 2912
rect 2814 2908 2818 2912
rect 2822 2898 2826 2902
rect 2694 2888 2698 2892
rect 2750 2888 2754 2892
rect 2726 2878 2730 2882
rect 2758 2878 2762 2882
rect 2782 2878 2786 2882
rect 2470 2868 2474 2872
rect 2486 2868 2490 2872
rect 2526 2868 2530 2872
rect 2574 2868 2578 2872
rect 2670 2868 2674 2872
rect 2686 2868 2690 2872
rect 2710 2868 2714 2872
rect 2494 2858 2498 2862
rect 2550 2858 2554 2862
rect 2598 2858 2602 2862
rect 2406 2838 2410 2842
rect 2366 2798 2370 2802
rect 2454 2848 2458 2852
rect 2470 2848 2474 2852
rect 2582 2848 2586 2852
rect 2438 2828 2442 2832
rect 2638 2858 2642 2862
rect 2702 2858 2706 2862
rect 2662 2848 2666 2852
rect 2686 2848 2690 2852
rect 2670 2838 2674 2842
rect 2614 2828 2618 2832
rect 2694 2818 2698 2822
rect 2486 2808 2490 2812
rect 2574 2808 2578 2812
rect 2538 2803 2542 2807
rect 2545 2803 2549 2807
rect 2446 2788 2450 2792
rect 2374 2778 2378 2782
rect 2422 2778 2426 2782
rect 2430 2778 2434 2782
rect 2342 2748 2346 2752
rect 2334 2738 2338 2742
rect 2326 2728 2330 2732
rect 2350 2728 2354 2732
rect 2318 2718 2322 2722
rect 2318 2668 2322 2672
rect 2230 2608 2234 2612
rect 2302 2608 2306 2612
rect 2262 2578 2266 2582
rect 2150 2568 2154 2572
rect 2174 2568 2178 2572
rect 2190 2548 2194 2552
rect 2166 2538 2170 2542
rect 2158 2528 2162 2532
rect 2190 2528 2194 2532
rect 2262 2558 2266 2562
rect 2286 2558 2290 2562
rect 2222 2548 2226 2552
rect 2278 2548 2282 2552
rect 2294 2548 2298 2552
rect 2214 2528 2218 2532
rect 2174 2518 2178 2522
rect 2198 2518 2202 2522
rect 2158 2508 2162 2512
rect 2206 2478 2210 2482
rect 2070 2468 2074 2472
rect 2230 2468 2234 2472
rect 2134 2448 2138 2452
rect 2190 2448 2194 2452
rect 2222 2448 2226 2452
rect 2086 2438 2090 2442
rect 2102 2438 2106 2442
rect 2134 2438 2138 2442
rect 2158 2438 2162 2442
rect 2182 2438 2186 2442
rect 1958 2418 1962 2422
rect 1886 2408 1890 2412
rect 1902 2408 1906 2412
rect 2070 2408 2074 2412
rect 1926 2388 1930 2392
rect 1774 2368 1778 2372
rect 1886 2368 1890 2372
rect 1910 2368 1914 2372
rect 2054 2368 2058 2372
rect 2070 2368 2074 2372
rect 2094 2368 2098 2372
rect 1718 2358 1722 2362
rect 1742 2358 1746 2362
rect 1798 2358 1802 2362
rect 1822 2348 1826 2352
rect 1718 2338 1722 2342
rect 1734 2338 1738 2342
rect 1750 2338 1754 2342
rect 1766 2338 1770 2342
rect 1782 2338 1786 2342
rect 1798 2338 1802 2342
rect 1758 2328 1762 2332
rect 1774 2328 1778 2332
rect 1790 2308 1794 2312
rect 1726 2298 1730 2302
rect 1750 2298 1754 2302
rect 1766 2298 1770 2302
rect 1718 2278 1722 2282
rect 1742 2278 1746 2282
rect 1686 2248 1690 2252
rect 1694 2248 1698 2252
rect 1678 2218 1682 2222
rect 1670 2178 1674 2182
rect 1662 2168 1666 2172
rect 1654 2158 1658 2162
rect 1614 2148 1618 2152
rect 1646 2148 1650 2152
rect 1574 2138 1578 2142
rect 1622 2138 1626 2142
rect 1638 2138 1642 2142
rect 1750 2248 1754 2252
rect 1782 2278 1786 2282
rect 1846 2328 1850 2332
rect 1870 2328 1874 2332
rect 1830 2308 1834 2312
rect 1830 2298 1834 2302
rect 1814 2288 1818 2292
rect 1798 2278 1802 2282
rect 1846 2288 1850 2292
rect 1838 2278 1842 2282
rect 1878 2278 1882 2282
rect 1862 2268 1866 2272
rect 1798 2248 1802 2252
rect 1822 2248 1826 2252
rect 1710 2208 1714 2212
rect 1718 2188 1722 2192
rect 1750 2188 1754 2192
rect 1702 2158 1706 2162
rect 1574 2118 1578 2122
rect 1582 2118 1586 2122
rect 1550 2098 1554 2102
rect 1606 2108 1610 2112
rect 1590 2078 1594 2082
rect 1630 2088 1634 2092
rect 1566 2068 1570 2072
rect 1606 2058 1610 2062
rect 1438 2038 1442 2042
rect 1502 2038 1506 2042
rect 1510 2038 1514 2042
rect 1406 2028 1410 2032
rect 1326 1958 1330 1962
rect 1334 1958 1338 1962
rect 1294 1948 1298 1952
rect 1246 1938 1250 1942
rect 1294 1928 1298 1932
rect 1310 1928 1314 1932
rect 1342 1948 1346 1952
rect 1358 1948 1362 1952
rect 1214 1908 1218 1912
rect 1222 1908 1226 1912
rect 1150 1878 1154 1882
rect 1166 1878 1170 1882
rect 1182 1878 1186 1882
rect 1174 1868 1178 1872
rect 1206 1868 1210 1872
rect 1126 1848 1130 1852
rect 1118 1788 1122 1792
rect 1110 1728 1114 1732
rect 1086 1708 1090 1712
rect 1102 1708 1106 1712
rect 1118 1708 1122 1712
rect 1102 1678 1106 1682
rect 1086 1668 1090 1672
rect 1286 1908 1290 1912
rect 1230 1888 1234 1892
rect 1230 1878 1234 1882
rect 1278 1878 1282 1882
rect 1254 1868 1258 1872
rect 1406 2008 1410 2012
rect 1374 1998 1378 2002
rect 1514 2003 1518 2007
rect 1521 2003 1525 2007
rect 1566 2048 1570 2052
rect 1638 2038 1642 2042
rect 1598 2028 1602 2032
rect 1478 1998 1482 2002
rect 1534 1998 1538 2002
rect 1462 1968 1466 1972
rect 1662 2118 1666 2122
rect 1686 2088 1690 2092
rect 1678 2058 1682 2062
rect 1734 2128 1738 2132
rect 1782 2198 1786 2202
rect 1798 2198 1802 2202
rect 1838 2198 1842 2202
rect 1766 2158 1770 2162
rect 1790 2178 1794 2182
rect 1830 2178 1834 2182
rect 1782 2138 1786 2142
rect 1814 2138 1818 2142
rect 1782 2128 1786 2132
rect 1758 2118 1762 2122
rect 1726 2098 1730 2102
rect 1718 2088 1722 2092
rect 1750 2108 1754 2112
rect 1694 2038 1698 2042
rect 1678 2028 1682 2032
rect 1646 2018 1650 2022
rect 1734 2018 1738 2022
rect 1542 1978 1546 1982
rect 1470 1958 1474 1962
rect 1518 1958 1522 1962
rect 1542 1958 1546 1962
rect 1382 1948 1386 1952
rect 1366 1928 1370 1932
rect 1382 1928 1386 1932
rect 1318 1888 1322 1892
rect 1318 1878 1322 1882
rect 1134 1838 1138 1842
rect 1214 1838 1218 1842
rect 1262 1848 1266 1852
rect 1294 1838 1298 1842
rect 1246 1828 1250 1832
rect 1222 1818 1226 1822
rect 1174 1798 1178 1802
rect 1190 1798 1194 1802
rect 1222 1798 1226 1802
rect 1134 1788 1138 1792
rect 1190 1788 1194 1792
rect 1158 1758 1162 1762
rect 1294 1798 1298 1802
rect 1286 1758 1290 1762
rect 1134 1738 1138 1742
rect 1134 1708 1138 1712
rect 1206 1748 1210 1752
rect 1270 1748 1274 1752
rect 1286 1748 1290 1752
rect 1182 1738 1186 1742
rect 1230 1738 1234 1742
rect 1278 1738 1282 1742
rect 1214 1728 1218 1732
rect 1270 1728 1274 1732
rect 1158 1718 1162 1722
rect 1190 1718 1194 1722
rect 1158 1698 1162 1702
rect 1150 1668 1154 1672
rect 1094 1658 1098 1662
rect 1126 1658 1130 1662
rect 1046 1648 1050 1652
rect 1022 1618 1026 1622
rect 1006 1608 1010 1612
rect 1046 1608 1050 1612
rect 1070 1608 1074 1612
rect 982 1568 986 1572
rect 1014 1598 1018 1602
rect 910 1478 914 1482
rect 918 1478 922 1482
rect 942 1478 946 1482
rect 950 1478 954 1482
rect 926 1468 930 1472
rect 902 1458 906 1462
rect 926 1448 930 1452
rect 726 1428 730 1432
rect 726 1348 730 1352
rect 750 1398 754 1402
rect 790 1398 794 1402
rect 718 1338 722 1342
rect 742 1318 746 1322
rect 702 1308 706 1312
rect 782 1368 786 1372
rect 878 1438 882 1442
rect 926 1438 930 1442
rect 838 1428 842 1432
rect 806 1388 810 1392
rect 798 1378 802 1382
rect 894 1378 898 1382
rect 958 1378 962 1382
rect 798 1368 802 1372
rect 838 1368 842 1372
rect 854 1368 858 1372
rect 878 1368 882 1372
rect 894 1368 898 1372
rect 758 1348 762 1352
rect 702 1298 706 1302
rect 710 1298 714 1302
rect 734 1298 738 1302
rect 750 1298 754 1302
rect 718 1268 722 1272
rect 694 1248 698 1252
rect 718 1248 722 1252
rect 686 1228 690 1232
rect 654 1178 658 1182
rect 742 1268 746 1272
rect 750 1198 754 1202
rect 734 1158 738 1162
rect 678 1148 682 1152
rect 694 1148 698 1152
rect 726 1148 730 1152
rect 822 1338 826 1342
rect 790 1278 794 1282
rect 806 1278 810 1282
rect 830 1328 834 1332
rect 846 1298 850 1302
rect 862 1338 866 1342
rect 782 1268 786 1272
rect 798 1268 802 1272
rect 822 1268 826 1272
rect 838 1268 842 1272
rect 806 1258 810 1262
rect 774 1228 778 1232
rect 798 1228 802 1232
rect 782 1208 786 1212
rect 774 1188 778 1192
rect 814 1188 818 1192
rect 766 1158 770 1162
rect 646 1138 650 1142
rect 654 1138 658 1142
rect 694 1138 698 1142
rect 742 1138 746 1142
rect 750 1138 754 1142
rect 758 1138 762 1142
rect 638 1098 642 1102
rect 638 1058 642 1062
rect 654 1058 658 1062
rect 686 1128 690 1132
rect 750 1128 754 1132
rect 734 1108 738 1112
rect 694 1098 698 1102
rect 686 1078 690 1082
rect 670 1068 674 1072
rect 662 1048 666 1052
rect 678 1048 682 1052
rect 662 1038 666 1042
rect 566 928 570 932
rect 614 928 618 932
rect 646 928 650 932
rect 558 898 562 902
rect 518 878 522 882
rect 534 878 538 882
rect 430 868 434 872
rect 470 868 474 872
rect 502 868 506 872
rect 358 808 362 812
rect 406 818 410 822
rect 422 808 426 812
rect 398 798 402 802
rect 454 838 458 842
rect 294 758 298 762
rect 366 758 370 762
rect 390 758 394 762
rect 422 758 426 762
rect 438 758 442 762
rect 254 738 258 742
rect 174 728 178 732
rect 182 728 186 732
rect 206 698 210 702
rect 278 748 282 752
rect 358 748 362 752
rect 390 748 394 752
rect 302 738 306 742
rect 270 718 274 722
rect 254 698 258 702
rect 182 678 186 682
rect 190 678 194 682
rect 302 728 306 732
rect 134 668 138 672
rect 198 668 202 672
rect 278 668 282 672
rect 62 638 66 642
rect 54 588 58 592
rect 46 548 50 552
rect 22 468 26 472
rect 30 468 34 472
rect 46 468 50 472
rect 22 458 26 462
rect 30 408 34 412
rect 22 378 26 382
rect 6 358 10 362
rect 70 558 74 562
rect 62 518 66 522
rect 86 628 90 632
rect 110 568 114 572
rect 102 558 106 562
rect 94 478 98 482
rect 94 468 98 472
rect 86 448 90 452
rect 142 658 146 662
rect 182 658 186 662
rect 150 628 154 632
rect 150 618 154 622
rect 142 608 146 612
rect 134 558 138 562
rect 118 498 122 502
rect 150 578 154 582
rect 182 598 186 602
rect 238 658 242 662
rect 214 638 218 642
rect 166 558 170 562
rect 166 478 170 482
rect 214 538 218 542
rect 198 528 202 532
rect 230 628 234 632
rect 254 648 258 652
rect 262 648 266 652
rect 270 588 274 592
rect 238 558 242 562
rect 206 478 210 482
rect 230 468 234 472
rect 166 448 170 452
rect 182 438 186 442
rect 206 428 210 432
rect 254 508 258 512
rect 262 488 266 492
rect 374 738 378 742
rect 318 678 322 682
rect 286 648 290 652
rect 294 648 298 652
rect 286 558 290 562
rect 310 558 314 562
rect 350 718 354 722
rect 366 678 370 682
rect 334 668 338 672
rect 342 658 346 662
rect 414 728 418 732
rect 414 678 418 682
rect 390 658 394 662
rect 382 638 386 642
rect 390 638 394 642
rect 374 608 378 612
rect 414 618 418 622
rect 334 578 338 582
rect 374 578 378 582
rect 430 728 434 732
rect 438 708 442 712
rect 510 848 514 852
rect 518 848 522 852
rect 494 838 498 842
rect 526 828 530 832
rect 482 803 486 807
rect 489 803 493 807
rect 470 798 474 802
rect 502 778 506 782
rect 462 748 466 752
rect 478 748 482 752
rect 518 748 522 752
rect 462 728 466 732
rect 462 718 466 722
rect 470 708 474 712
rect 454 658 458 662
rect 462 658 466 662
rect 430 638 434 642
rect 430 628 434 632
rect 422 568 426 572
rect 334 558 338 562
rect 318 538 322 542
rect 294 518 298 522
rect 326 488 330 492
rect 302 478 306 482
rect 358 528 362 532
rect 366 518 370 522
rect 334 478 338 482
rect 502 688 506 692
rect 486 678 490 682
rect 606 918 610 922
rect 718 1068 722 1072
rect 718 1058 722 1062
rect 694 1018 698 1022
rect 710 1018 714 1022
rect 678 1008 682 1012
rect 798 1158 802 1162
rect 838 1258 842 1262
rect 806 1148 810 1152
rect 822 1148 826 1152
rect 878 1328 882 1332
rect 994 1503 998 1507
rect 1001 1503 1005 1507
rect 974 1478 978 1482
rect 982 1478 986 1482
rect 1038 1588 1042 1592
rect 1030 1548 1034 1552
rect 1078 1578 1082 1582
rect 1094 1578 1098 1582
rect 1070 1568 1074 1572
rect 1086 1568 1090 1572
rect 1086 1548 1090 1552
rect 1102 1548 1106 1552
rect 1022 1538 1026 1542
rect 1046 1538 1050 1542
rect 1062 1538 1066 1542
rect 1094 1538 1098 1542
rect 1086 1518 1090 1522
rect 1022 1508 1026 1512
rect 1030 1488 1034 1492
rect 1030 1478 1034 1482
rect 998 1458 1002 1462
rect 1006 1458 1010 1462
rect 1022 1458 1026 1462
rect 974 1428 978 1432
rect 974 1388 978 1392
rect 1022 1428 1026 1432
rect 1014 1398 1018 1402
rect 926 1358 930 1362
rect 966 1358 970 1362
rect 990 1358 994 1362
rect 998 1358 1002 1362
rect 902 1348 906 1352
rect 974 1348 978 1352
rect 1006 1348 1010 1352
rect 1014 1348 1018 1352
rect 910 1338 914 1342
rect 950 1338 954 1342
rect 878 1308 882 1312
rect 894 1278 898 1282
rect 854 1258 858 1262
rect 870 1258 874 1262
rect 870 1198 874 1202
rect 846 1158 850 1162
rect 798 1138 802 1142
rect 814 1138 818 1142
rect 846 1138 850 1142
rect 774 1128 778 1132
rect 790 1128 794 1132
rect 774 1118 778 1122
rect 830 1118 834 1122
rect 822 1088 826 1092
rect 742 1068 746 1072
rect 758 1068 762 1072
rect 750 1058 754 1062
rect 742 1018 746 1022
rect 710 998 714 1002
rect 734 998 738 1002
rect 686 988 690 992
rect 670 908 674 912
rect 598 888 602 892
rect 630 888 634 892
rect 582 868 586 872
rect 550 858 554 862
rect 566 768 570 772
rect 630 878 634 882
rect 614 868 618 872
rect 630 858 634 862
rect 622 848 626 852
rect 582 838 586 842
rect 598 838 602 842
rect 614 838 618 842
rect 598 818 602 822
rect 614 818 618 822
rect 582 768 586 772
rect 550 748 554 752
rect 574 748 578 752
rect 542 738 546 742
rect 526 678 530 682
rect 542 678 546 682
rect 558 738 562 742
rect 566 738 570 742
rect 582 738 586 742
rect 558 658 562 662
rect 518 648 522 652
rect 510 638 514 642
rect 534 638 538 642
rect 478 628 482 632
rect 482 603 486 607
rect 489 603 493 607
rect 502 558 506 562
rect 542 558 546 562
rect 518 548 522 552
rect 414 538 418 542
rect 414 528 418 532
rect 422 528 426 532
rect 390 518 394 522
rect 382 508 386 512
rect 414 508 418 512
rect 406 478 410 482
rect 278 468 282 472
rect 286 468 290 472
rect 358 468 362 472
rect 390 468 394 472
rect 302 458 306 462
rect 366 458 370 462
rect 382 458 386 462
rect 398 458 402 462
rect 414 458 418 462
rect 246 438 250 442
rect 230 418 234 422
rect 222 408 226 412
rect 102 358 106 362
rect 38 348 42 352
rect 62 348 66 352
rect 134 348 138 352
rect 174 348 178 352
rect 182 348 186 352
rect 86 288 90 292
rect 158 338 162 342
rect 190 338 194 342
rect 238 388 242 392
rect 182 328 186 332
rect 206 328 210 332
rect 174 318 178 322
rect 166 268 170 272
rect 62 258 66 262
rect 6 248 10 252
rect 30 248 34 252
rect 70 248 74 252
rect 54 178 58 182
rect 110 238 114 242
rect 110 178 114 182
rect 214 288 218 292
rect 246 328 250 332
rect 310 438 314 442
rect 342 438 346 442
rect 278 418 282 422
rect 334 408 338 412
rect 366 398 370 402
rect 262 358 266 362
rect 278 338 282 342
rect 294 298 298 302
rect 214 268 218 272
rect 182 228 186 232
rect 182 218 186 222
rect 150 198 154 202
rect 30 148 34 152
rect 30 68 34 72
rect 54 88 58 92
rect 102 138 106 142
rect 134 138 138 142
rect 166 138 170 142
rect 198 138 202 142
rect 118 88 122 92
rect 214 128 218 132
rect 158 88 162 92
rect 6 58 10 62
rect 46 58 50 62
rect 206 58 210 62
rect 70 48 74 52
rect 102 48 106 52
rect 86 28 90 32
rect 262 238 266 242
rect 318 338 322 342
rect 334 338 338 342
rect 350 338 354 342
rect 350 318 354 322
rect 382 338 386 342
rect 366 328 370 332
rect 374 328 378 332
rect 310 268 314 272
rect 358 268 362 272
rect 390 318 394 322
rect 374 268 378 272
rect 286 248 290 252
rect 318 248 322 252
rect 278 238 282 242
rect 270 218 274 222
rect 318 208 322 212
rect 310 168 314 172
rect 302 158 306 162
rect 246 108 250 112
rect 222 48 226 52
rect 246 48 250 52
rect 278 138 282 142
rect 286 128 290 132
rect 270 98 274 102
rect 278 98 282 102
rect 326 178 330 182
rect 334 158 338 162
rect 406 268 410 272
rect 430 428 434 432
rect 470 518 474 522
rect 454 508 458 512
rect 462 428 466 432
rect 454 418 458 422
rect 558 608 562 612
rect 638 828 642 832
rect 630 798 634 802
rect 646 748 650 752
rect 622 738 626 742
rect 606 688 610 692
rect 622 698 626 702
rect 590 658 594 662
rect 606 658 610 662
rect 582 628 586 632
rect 582 578 586 582
rect 550 518 554 522
rect 614 638 618 642
rect 614 618 618 622
rect 638 718 642 722
rect 694 978 698 982
rect 694 948 698 952
rect 702 878 706 882
rect 686 848 690 852
rect 678 838 682 842
rect 662 828 666 832
rect 678 788 682 792
rect 782 1068 786 1072
rect 806 1068 810 1072
rect 790 1058 794 1062
rect 758 1028 762 1032
rect 774 1028 778 1032
rect 726 938 730 942
rect 806 1048 810 1052
rect 814 1048 818 1052
rect 886 1158 890 1162
rect 878 1138 882 1142
rect 886 1128 890 1132
rect 862 1118 866 1122
rect 854 1108 858 1112
rect 878 1088 882 1092
rect 830 1068 834 1072
rect 846 1068 850 1072
rect 926 1298 930 1302
rect 982 1338 986 1342
rect 982 1308 986 1312
rect 974 1298 978 1302
rect 934 1278 938 1282
rect 966 1278 970 1282
rect 974 1278 978 1282
rect 918 1258 922 1262
rect 902 1238 906 1242
rect 902 1218 906 1222
rect 966 1268 970 1272
rect 994 1303 998 1307
rect 1001 1303 1005 1307
rect 1014 1298 1018 1302
rect 982 1268 986 1272
rect 1054 1468 1058 1472
rect 1070 1478 1074 1482
rect 1134 1568 1138 1572
rect 1150 1628 1154 1632
rect 1150 1598 1154 1602
rect 1142 1528 1146 1532
rect 1126 1518 1130 1522
rect 1134 1518 1138 1522
rect 1118 1498 1122 1502
rect 1134 1498 1138 1502
rect 1230 1698 1234 1702
rect 1174 1668 1178 1672
rect 1214 1668 1218 1672
rect 1222 1668 1226 1672
rect 1342 1838 1346 1842
rect 1334 1828 1338 1832
rect 1358 1908 1362 1912
rect 1414 1948 1418 1952
rect 1422 1948 1426 1952
rect 1558 1948 1562 1952
rect 1446 1938 1450 1942
rect 1462 1928 1466 1932
rect 1430 1908 1434 1912
rect 1390 1888 1394 1892
rect 1430 1878 1434 1882
rect 1366 1868 1370 1872
rect 1374 1858 1378 1862
rect 1366 1808 1370 1812
rect 1350 1768 1354 1772
rect 1358 1768 1362 1772
rect 1342 1758 1346 1762
rect 1366 1758 1370 1762
rect 1302 1748 1306 1752
rect 1326 1738 1330 1742
rect 1318 1728 1322 1732
rect 1302 1718 1306 1722
rect 1262 1668 1266 1672
rect 1198 1658 1202 1662
rect 1270 1658 1274 1662
rect 1174 1598 1178 1602
rect 1158 1528 1162 1532
rect 1174 1528 1178 1532
rect 1174 1518 1178 1522
rect 1166 1508 1170 1512
rect 1278 1648 1282 1652
rect 1286 1648 1290 1652
rect 1254 1618 1258 1622
rect 1262 1618 1266 1622
rect 1238 1608 1242 1612
rect 1222 1598 1226 1602
rect 1246 1598 1250 1602
rect 1230 1588 1234 1592
rect 1262 1588 1266 1592
rect 1326 1698 1330 1702
rect 1326 1678 1330 1682
rect 1342 1678 1346 1682
rect 1446 1868 1450 1872
rect 1422 1858 1426 1862
rect 1390 1838 1394 1842
rect 1462 1848 1466 1852
rect 1438 1828 1442 1832
rect 1422 1818 1426 1822
rect 1454 1818 1458 1822
rect 1398 1808 1402 1812
rect 1382 1778 1386 1782
rect 1390 1758 1394 1762
rect 1366 1738 1370 1742
rect 1382 1738 1386 1742
rect 1446 1808 1450 1812
rect 1462 1808 1466 1812
rect 1446 1758 1450 1762
rect 1406 1748 1410 1752
rect 1414 1748 1418 1752
rect 1398 1738 1402 1742
rect 1318 1668 1322 1672
rect 1374 1678 1378 1682
rect 1390 1668 1394 1672
rect 1422 1728 1426 1732
rect 1406 1708 1410 1712
rect 1494 1938 1498 1942
rect 1542 1938 1546 1942
rect 1558 1938 1562 1942
rect 1566 1938 1570 1942
rect 1582 1938 1586 1942
rect 1542 1928 1546 1932
rect 1550 1928 1554 1932
rect 1574 1928 1578 1932
rect 1502 1908 1506 1912
rect 1494 1888 1498 1892
rect 1550 1888 1554 1892
rect 1486 1868 1490 1872
rect 1486 1858 1490 1862
rect 1518 1858 1522 1862
rect 1534 1858 1538 1862
rect 1502 1838 1506 1842
rect 1486 1738 1490 1742
rect 1454 1718 1458 1722
rect 1438 1708 1442 1712
rect 1478 1698 1482 1702
rect 1430 1688 1434 1692
rect 1414 1668 1418 1672
rect 1334 1658 1338 1662
rect 1358 1658 1362 1662
rect 1406 1658 1410 1662
rect 1326 1648 1330 1652
rect 1350 1628 1354 1632
rect 1358 1628 1362 1632
rect 1334 1618 1338 1622
rect 1206 1568 1210 1572
rect 1222 1568 1226 1572
rect 1206 1548 1210 1552
rect 1246 1548 1250 1552
rect 1230 1538 1234 1542
rect 1198 1508 1202 1512
rect 1190 1488 1194 1492
rect 1126 1458 1130 1462
rect 1134 1458 1138 1462
rect 1158 1458 1162 1462
rect 1166 1458 1170 1462
rect 1030 1418 1034 1422
rect 1070 1448 1074 1452
rect 1094 1448 1098 1452
rect 1062 1378 1066 1382
rect 1062 1358 1066 1362
rect 1038 1338 1042 1342
rect 1054 1328 1058 1332
rect 1038 1288 1042 1292
rect 1054 1288 1058 1292
rect 1006 1268 1010 1272
rect 1014 1268 1018 1272
rect 1038 1268 1042 1272
rect 950 1258 954 1262
rect 982 1238 986 1242
rect 934 1198 938 1202
rect 950 1198 954 1202
rect 934 1188 938 1192
rect 950 1188 954 1192
rect 910 1138 914 1142
rect 918 1138 922 1142
rect 910 1118 914 1122
rect 894 1088 898 1092
rect 798 1018 802 1022
rect 822 1008 826 1012
rect 814 978 818 982
rect 798 958 802 962
rect 758 948 762 952
rect 782 948 786 952
rect 806 948 810 952
rect 718 878 722 882
rect 750 938 754 942
rect 782 938 786 942
rect 790 928 794 932
rect 742 868 746 872
rect 774 868 778 872
rect 726 858 730 862
rect 726 838 730 842
rect 750 838 754 842
rect 766 828 770 832
rect 774 828 778 832
rect 838 1058 842 1062
rect 862 1048 866 1052
rect 878 1048 882 1052
rect 854 948 858 952
rect 854 938 858 942
rect 966 1148 970 1152
rect 966 1138 970 1142
rect 942 1128 946 1132
rect 926 1118 930 1122
rect 942 1118 946 1122
rect 926 1098 930 1102
rect 1022 1258 1026 1262
rect 998 1198 1002 1202
rect 990 1188 994 1192
rect 1022 1238 1026 1242
rect 1038 1198 1042 1202
rect 1014 1148 1018 1152
rect 1022 1138 1026 1142
rect 1038 1138 1042 1142
rect 974 1118 978 1122
rect 950 1108 954 1112
rect 950 1088 954 1092
rect 918 1048 922 1052
rect 926 1048 930 1052
rect 886 1028 890 1032
rect 894 1018 898 1022
rect 894 1008 898 1012
rect 902 1008 906 1012
rect 878 948 882 952
rect 870 928 874 932
rect 830 918 834 922
rect 878 918 882 922
rect 798 898 802 902
rect 806 888 810 892
rect 822 888 826 892
rect 806 878 810 882
rect 798 858 802 862
rect 814 848 818 852
rect 838 888 842 892
rect 878 888 882 892
rect 830 878 834 882
rect 830 858 834 862
rect 854 858 858 862
rect 878 858 882 862
rect 846 838 850 842
rect 822 828 826 832
rect 846 828 850 832
rect 790 808 794 812
rect 806 808 810 812
rect 726 798 730 802
rect 782 798 786 802
rect 814 798 818 802
rect 742 778 746 782
rect 782 778 786 782
rect 718 768 722 772
rect 758 768 762 772
rect 670 738 674 742
rect 702 738 706 742
rect 742 738 746 742
rect 662 728 666 732
rect 694 728 698 732
rect 734 728 738 732
rect 718 698 722 702
rect 726 688 730 692
rect 750 688 754 692
rect 662 668 666 672
rect 678 668 682 672
rect 814 768 818 772
rect 822 758 826 762
rect 854 758 858 762
rect 846 748 850 752
rect 886 808 890 812
rect 886 798 890 802
rect 878 768 882 772
rect 902 998 906 1002
rect 910 988 914 992
rect 942 1048 946 1052
rect 950 1028 954 1032
rect 934 1018 938 1022
rect 942 998 946 1002
rect 966 1078 970 1082
rect 994 1103 998 1107
rect 1001 1103 1005 1107
rect 1030 1128 1034 1132
rect 1022 1108 1026 1112
rect 1014 1088 1018 1092
rect 982 1068 986 1072
rect 990 1058 994 1062
rect 1022 1058 1026 1062
rect 966 1018 970 1022
rect 974 1018 978 1022
rect 1014 1018 1018 1022
rect 958 998 962 1002
rect 966 998 970 1002
rect 1014 998 1018 1002
rect 966 988 970 992
rect 1014 978 1018 982
rect 918 948 922 952
rect 950 948 954 952
rect 910 928 914 932
rect 950 908 954 912
rect 966 908 970 912
rect 926 898 930 902
rect 942 898 946 902
rect 982 948 986 952
rect 990 938 994 942
rect 982 908 986 912
rect 918 888 922 892
rect 934 888 938 892
rect 910 878 914 882
rect 958 878 962 882
rect 950 868 954 872
rect 918 838 922 842
rect 950 838 954 842
rect 926 828 930 832
rect 902 808 906 812
rect 918 768 922 772
rect 926 768 930 772
rect 934 768 938 772
rect 894 758 898 762
rect 902 758 906 762
rect 974 858 978 862
rect 966 838 970 842
rect 994 903 998 907
rect 1001 903 1005 907
rect 998 888 1002 892
rect 1078 1428 1082 1432
rect 1110 1428 1114 1432
rect 1086 1418 1090 1422
rect 1094 1348 1098 1352
rect 1118 1418 1122 1422
rect 1102 1328 1106 1332
rect 1158 1438 1162 1442
rect 1174 1438 1178 1442
rect 1166 1388 1170 1392
rect 1134 1358 1138 1362
rect 1158 1358 1162 1362
rect 1070 1278 1074 1282
rect 1094 1278 1098 1282
rect 1062 1268 1066 1272
rect 1102 1268 1106 1272
rect 1070 1258 1074 1262
rect 1094 1258 1098 1262
rect 1094 1228 1098 1232
rect 1054 1198 1058 1202
rect 1062 1198 1066 1202
rect 1054 1148 1058 1152
rect 1078 1198 1082 1202
rect 1078 1138 1082 1142
rect 1078 1098 1082 1102
rect 1102 1178 1106 1182
rect 1086 1088 1090 1092
rect 1038 1058 1042 1062
rect 1046 1058 1050 1062
rect 1038 1008 1042 1012
rect 1046 998 1050 1002
rect 1086 1068 1090 1072
rect 1150 1338 1154 1342
rect 1134 1308 1138 1312
rect 1126 1298 1130 1302
rect 1198 1448 1202 1452
rect 1190 1418 1194 1422
rect 1190 1368 1194 1372
rect 1222 1488 1226 1492
rect 1214 1468 1218 1472
rect 1278 1578 1282 1582
rect 1302 1588 1306 1592
rect 1318 1588 1322 1592
rect 1334 1558 1338 1562
rect 1318 1548 1322 1552
rect 1326 1548 1330 1552
rect 1302 1538 1306 1542
rect 1254 1528 1258 1532
rect 1262 1528 1266 1532
rect 1286 1528 1290 1532
rect 1294 1528 1298 1532
rect 1310 1528 1314 1532
rect 1302 1518 1306 1522
rect 1262 1478 1266 1482
rect 1278 1478 1282 1482
rect 1302 1488 1306 1492
rect 1302 1478 1306 1482
rect 1286 1468 1290 1472
rect 1222 1458 1226 1462
rect 1246 1458 1250 1462
rect 1310 1458 1314 1462
rect 1278 1438 1282 1442
rect 1254 1418 1258 1422
rect 1270 1398 1274 1402
rect 1278 1398 1282 1402
rect 1310 1398 1314 1402
rect 1238 1378 1242 1382
rect 1262 1378 1266 1382
rect 1206 1348 1210 1352
rect 1238 1348 1242 1352
rect 1182 1328 1186 1332
rect 1198 1328 1202 1332
rect 1214 1328 1218 1332
rect 1222 1328 1226 1332
rect 1158 1288 1162 1292
rect 1190 1298 1194 1302
rect 1166 1278 1170 1282
rect 1126 1268 1130 1272
rect 1158 1268 1162 1272
rect 1142 1248 1146 1252
rect 1126 1188 1130 1192
rect 1126 1168 1130 1172
rect 1158 1258 1162 1262
rect 1174 1258 1178 1262
rect 1166 1248 1170 1252
rect 1166 1218 1170 1222
rect 1158 1178 1162 1182
rect 1142 1148 1146 1152
rect 1118 1108 1122 1112
rect 1118 1088 1122 1092
rect 1110 1078 1114 1082
rect 1110 1068 1114 1072
rect 1126 1068 1130 1072
rect 1062 1058 1066 1062
rect 1102 1058 1106 1062
rect 1070 1048 1074 1052
rect 1206 1288 1210 1292
rect 1222 1278 1226 1282
rect 1222 1268 1226 1272
rect 1214 1258 1218 1262
rect 1214 1238 1218 1242
rect 1190 1228 1194 1232
rect 1222 1228 1226 1232
rect 1198 1218 1202 1222
rect 1214 1218 1218 1222
rect 1182 1188 1186 1192
rect 1174 1178 1178 1182
rect 1214 1178 1218 1182
rect 1206 1168 1210 1172
rect 1174 1158 1178 1162
rect 1182 1138 1186 1142
rect 1166 1128 1170 1132
rect 1190 1128 1194 1132
rect 1142 1088 1146 1092
rect 1174 1058 1178 1062
rect 1158 1048 1162 1052
rect 1110 1038 1114 1042
rect 1102 1008 1106 1012
rect 1054 988 1058 992
rect 1086 988 1090 992
rect 1038 978 1042 982
rect 1078 978 1082 982
rect 1062 968 1066 972
rect 1030 928 1034 932
rect 1022 908 1026 912
rect 1046 938 1050 942
rect 1206 1138 1210 1142
rect 1214 1108 1218 1112
rect 1270 1358 1274 1362
rect 1286 1358 1290 1362
rect 1302 1358 1306 1362
rect 1310 1338 1314 1342
rect 1270 1318 1274 1322
rect 1278 1318 1282 1322
rect 1262 1288 1266 1292
rect 1278 1288 1282 1292
rect 1302 1288 1306 1292
rect 1254 1278 1258 1282
rect 1390 1628 1394 1632
rect 1374 1618 1378 1622
rect 1366 1598 1370 1602
rect 1366 1548 1370 1552
rect 1350 1528 1354 1532
rect 1342 1498 1346 1502
rect 1342 1478 1346 1482
rect 1398 1598 1402 1602
rect 1514 1803 1518 1807
rect 1521 1803 1525 1807
rect 1510 1778 1514 1782
rect 1542 1818 1546 1822
rect 1566 1818 1570 1822
rect 1534 1768 1538 1772
rect 1518 1748 1522 1752
rect 1526 1728 1530 1732
rect 1558 1728 1562 1732
rect 1566 1718 1570 1722
rect 1550 1708 1554 1712
rect 1550 1698 1554 1702
rect 1590 1928 1594 1932
rect 1598 1928 1602 1932
rect 1630 1998 1634 2002
rect 1622 1958 1626 1962
rect 1614 1898 1618 1902
rect 1678 2008 1682 2012
rect 1694 2008 1698 2012
rect 1678 1978 1682 1982
rect 1654 1958 1658 1962
rect 1662 1948 1666 1952
rect 1646 1938 1650 1942
rect 1638 1928 1642 1932
rect 1638 1878 1642 1882
rect 1686 1968 1690 1972
rect 1694 1958 1698 1962
rect 1806 2098 1810 2102
rect 1814 2098 1818 2102
rect 1782 2068 1786 2072
rect 1726 1978 1730 1982
rect 1718 1968 1722 1972
rect 1742 1968 1746 1972
rect 1750 1968 1754 1972
rect 1726 1958 1730 1962
rect 1686 1938 1690 1942
rect 1662 1898 1666 1902
rect 1678 1898 1682 1902
rect 1582 1868 1586 1872
rect 1646 1868 1650 1872
rect 1598 1858 1602 1862
rect 1590 1848 1594 1852
rect 1614 1848 1618 1852
rect 1622 1848 1626 1852
rect 1638 1828 1642 1832
rect 1598 1808 1602 1812
rect 1606 1808 1610 1812
rect 1646 1808 1650 1812
rect 1670 1858 1674 1862
rect 1670 1848 1674 1852
rect 1670 1828 1674 1832
rect 1718 1938 1722 1942
rect 1710 1908 1714 1912
rect 1702 1898 1706 1902
rect 1774 2048 1778 2052
rect 1974 2358 1978 2362
rect 1894 2348 1898 2352
rect 1934 2348 1938 2352
rect 1974 2348 1978 2352
rect 1982 2348 1986 2352
rect 2030 2348 2034 2352
rect 2046 2348 2050 2352
rect 1918 2338 1922 2342
rect 1950 2338 1954 2342
rect 1902 2328 1906 2332
rect 1998 2338 2002 2342
rect 1942 2308 1946 2312
rect 2006 2318 2010 2322
rect 1998 2308 2002 2312
rect 1902 2278 1906 2282
rect 1958 2278 1962 2282
rect 1974 2278 1978 2282
rect 1878 2198 1882 2202
rect 1902 2268 1906 2272
rect 1942 2258 1946 2262
rect 2026 2303 2030 2307
rect 2033 2303 2037 2307
rect 2046 2298 2050 2302
rect 2014 2278 2018 2282
rect 2150 2398 2154 2402
rect 2110 2358 2114 2362
rect 2070 2328 2074 2332
rect 2086 2328 2090 2332
rect 2102 2328 2106 2332
rect 2110 2328 2114 2332
rect 2134 2328 2138 2332
rect 2078 2308 2082 2312
rect 2030 2258 2034 2262
rect 1966 2248 1970 2252
rect 1910 2198 1914 2202
rect 1966 2198 1970 2202
rect 1886 2168 1890 2172
rect 1870 2158 1874 2162
rect 1854 2148 1858 2152
rect 1950 2168 1954 2172
rect 1918 2158 1922 2162
rect 1966 2158 1970 2162
rect 2078 2268 2082 2272
rect 2014 2198 2018 2202
rect 2142 2318 2146 2322
rect 2158 2358 2162 2362
rect 2238 2448 2242 2452
rect 2238 2438 2242 2442
rect 2214 2408 2218 2412
rect 2198 2388 2202 2392
rect 2190 2358 2194 2362
rect 2198 2348 2202 2352
rect 2166 2338 2170 2342
rect 2182 2308 2186 2312
rect 2262 2528 2266 2532
rect 2286 2518 2290 2522
rect 2254 2498 2258 2502
rect 2254 2468 2258 2472
rect 2270 2448 2274 2452
rect 2262 2438 2266 2442
rect 2246 2418 2250 2422
rect 2326 2578 2330 2582
rect 2310 2568 2314 2572
rect 2414 2758 2418 2762
rect 2382 2748 2386 2752
rect 2566 2778 2570 2782
rect 2502 2768 2506 2772
rect 2446 2758 2450 2762
rect 2462 2758 2466 2762
rect 2526 2758 2530 2762
rect 2558 2758 2562 2762
rect 2438 2718 2442 2722
rect 2430 2708 2434 2712
rect 2358 2698 2362 2702
rect 2454 2748 2458 2752
rect 2510 2748 2514 2752
rect 2462 2738 2466 2742
rect 2502 2738 2506 2742
rect 2382 2688 2386 2692
rect 2398 2688 2402 2692
rect 2350 2678 2354 2682
rect 2366 2678 2370 2682
rect 2550 2698 2554 2702
rect 2342 2668 2346 2672
rect 2350 2618 2354 2622
rect 2398 2668 2402 2672
rect 2422 2666 2426 2670
rect 2382 2638 2386 2642
rect 2430 2618 2434 2622
rect 2406 2598 2410 2602
rect 2334 2558 2338 2562
rect 2342 2558 2346 2562
rect 2350 2558 2354 2562
rect 2462 2668 2466 2672
rect 2494 2668 2498 2672
rect 2502 2668 2506 2672
rect 2534 2668 2538 2672
rect 2558 2668 2562 2672
rect 2518 2658 2522 2662
rect 2470 2638 2474 2642
rect 2526 2638 2530 2642
rect 2518 2618 2522 2622
rect 2438 2568 2442 2572
rect 2454 2558 2458 2562
rect 2486 2558 2490 2562
rect 2502 2558 2506 2562
rect 2350 2538 2354 2542
rect 2398 2528 2402 2532
rect 2406 2528 2410 2532
rect 2374 2508 2378 2512
rect 2390 2508 2394 2512
rect 2398 2508 2402 2512
rect 2326 2488 2330 2492
rect 2342 2488 2346 2492
rect 2438 2548 2442 2552
rect 2438 2518 2442 2522
rect 2318 2468 2322 2472
rect 2342 2468 2346 2472
rect 2406 2468 2410 2472
rect 2438 2468 2442 2472
rect 2286 2438 2290 2442
rect 2294 2438 2298 2442
rect 2326 2448 2330 2452
rect 2358 2448 2362 2452
rect 2366 2448 2370 2452
rect 2318 2408 2322 2412
rect 2350 2438 2354 2442
rect 2374 2438 2378 2442
rect 2374 2408 2378 2412
rect 2390 2408 2394 2412
rect 2382 2398 2386 2402
rect 2538 2603 2542 2607
rect 2545 2603 2549 2607
rect 2526 2598 2530 2602
rect 2574 2738 2578 2742
rect 2582 2678 2586 2682
rect 2574 2668 2578 2672
rect 2566 2658 2570 2662
rect 2582 2658 2586 2662
rect 2574 2638 2578 2642
rect 2686 2778 2690 2782
rect 2598 2768 2602 2772
rect 2670 2758 2674 2762
rect 2662 2748 2666 2752
rect 2614 2728 2618 2732
rect 2638 2738 2642 2742
rect 2630 2718 2634 2722
rect 2670 2718 2674 2722
rect 2598 2708 2602 2712
rect 2662 2708 2666 2712
rect 2598 2698 2602 2702
rect 2614 2698 2618 2702
rect 2646 2698 2650 2702
rect 2654 2698 2658 2702
rect 2638 2688 2642 2692
rect 2678 2678 2682 2682
rect 2638 2668 2642 2672
rect 2606 2658 2610 2662
rect 2622 2658 2626 2662
rect 2630 2658 2634 2662
rect 2598 2608 2602 2612
rect 2590 2578 2594 2582
rect 2614 2578 2618 2582
rect 2558 2568 2562 2572
rect 2478 2538 2482 2542
rect 2494 2538 2498 2542
rect 2478 2518 2482 2522
rect 2518 2528 2522 2532
rect 2526 2528 2530 2532
rect 2470 2508 2474 2512
rect 2510 2508 2514 2512
rect 2462 2498 2466 2502
rect 2454 2488 2458 2492
rect 2454 2468 2458 2472
rect 2446 2458 2450 2462
rect 2414 2428 2418 2432
rect 2438 2428 2442 2432
rect 2326 2388 2330 2392
rect 2390 2388 2394 2392
rect 2414 2388 2418 2392
rect 2238 2368 2242 2372
rect 2270 2368 2274 2372
rect 2278 2368 2282 2372
rect 2222 2348 2226 2352
rect 2158 2288 2162 2292
rect 2198 2288 2202 2292
rect 2126 2278 2130 2282
rect 2142 2278 2146 2282
rect 2182 2278 2186 2282
rect 2110 2268 2114 2272
rect 2134 2268 2138 2272
rect 2062 2208 2066 2212
rect 2110 2208 2114 2212
rect 2118 2208 2122 2212
rect 2078 2198 2082 2202
rect 2030 2168 2034 2172
rect 2046 2168 2050 2172
rect 2006 2158 2010 2162
rect 1990 2148 1994 2152
rect 1846 2138 1850 2142
rect 1862 2138 1866 2142
rect 1918 2138 1922 2142
rect 1966 2138 1970 2142
rect 1982 2138 1986 2142
rect 1870 2118 1874 2122
rect 1974 2118 1978 2122
rect 2014 2118 2018 2122
rect 1862 2098 1866 2102
rect 1846 2058 1850 2062
rect 1822 2028 1826 2032
rect 1782 2018 1786 2022
rect 1782 1998 1786 2002
rect 1790 1998 1794 2002
rect 1766 1928 1770 1932
rect 1782 1928 1786 1932
rect 1758 1918 1762 1922
rect 1774 1918 1778 1922
rect 1782 1908 1786 1912
rect 1862 2048 1866 2052
rect 1886 2098 1890 2102
rect 1926 2098 1930 2102
rect 1878 2078 1882 2082
rect 1926 2078 1930 2082
rect 1958 2108 1962 2112
rect 2026 2103 2030 2107
rect 2033 2103 2037 2107
rect 1942 2068 1946 2072
rect 1998 2068 2002 2072
rect 2006 2068 2010 2072
rect 2014 2068 2018 2072
rect 1886 2058 1890 2062
rect 1902 2048 1906 2052
rect 1910 2048 1914 2052
rect 1854 2038 1858 2042
rect 1910 2018 1914 2022
rect 1870 2008 1874 2012
rect 1942 2048 1946 2052
rect 1982 2038 1986 2042
rect 2038 2038 2042 2042
rect 1950 2018 1954 2022
rect 1966 2018 1970 2022
rect 1934 2008 1938 2012
rect 1966 2008 1970 2012
rect 1950 1998 1954 2002
rect 1830 1978 1834 1982
rect 1846 1978 1850 1982
rect 1878 1978 1882 1982
rect 1958 1978 1962 1982
rect 1838 1958 1842 1962
rect 1862 1958 1866 1962
rect 1934 1958 1938 1962
rect 1950 1958 1954 1962
rect 1838 1948 1842 1952
rect 1846 1948 1850 1952
rect 1862 1948 1866 1952
rect 1942 1948 1946 1952
rect 1798 1928 1802 1932
rect 1822 1928 1826 1932
rect 1814 1918 1818 1922
rect 1822 1908 1826 1912
rect 1998 1948 2002 1952
rect 1966 1938 1970 1942
rect 1974 1938 1978 1942
rect 1878 1928 1882 1932
rect 1894 1928 1898 1932
rect 1902 1928 1906 1932
rect 1926 1928 1930 1932
rect 1870 1918 1874 1922
rect 1910 1918 1914 1922
rect 1942 1918 1946 1922
rect 1982 1918 1986 1922
rect 1838 1908 1842 1912
rect 1846 1908 1850 1912
rect 1854 1908 1858 1912
rect 1798 1898 1802 1902
rect 1806 1898 1810 1902
rect 1822 1898 1826 1902
rect 1830 1898 1834 1902
rect 1694 1858 1698 1862
rect 1710 1858 1714 1862
rect 1726 1858 1730 1862
rect 1750 1858 1754 1862
rect 1710 1848 1714 1852
rect 1686 1808 1690 1812
rect 1678 1798 1682 1802
rect 1654 1788 1658 1792
rect 1654 1768 1658 1772
rect 1590 1758 1594 1762
rect 1622 1758 1626 1762
rect 1638 1758 1642 1762
rect 1646 1758 1650 1762
rect 1590 1748 1594 1752
rect 1630 1748 1634 1752
rect 1582 1738 1586 1742
rect 1606 1738 1610 1742
rect 1638 1738 1642 1742
rect 1598 1728 1602 1732
rect 1638 1728 1642 1732
rect 1630 1698 1634 1702
rect 1598 1688 1602 1692
rect 1550 1678 1554 1682
rect 1430 1668 1434 1672
rect 1446 1668 1450 1672
rect 1494 1668 1498 1672
rect 1470 1658 1474 1662
rect 1566 1658 1570 1662
rect 1422 1628 1426 1632
rect 1438 1628 1442 1632
rect 1454 1628 1458 1632
rect 1478 1628 1482 1632
rect 1430 1598 1434 1602
rect 1390 1588 1394 1592
rect 1414 1588 1418 1592
rect 1406 1558 1410 1562
rect 1422 1558 1426 1562
rect 1382 1538 1386 1542
rect 1358 1478 1362 1482
rect 1406 1538 1410 1542
rect 1422 1538 1426 1542
rect 1398 1528 1402 1532
rect 1398 1518 1402 1522
rect 1390 1488 1394 1492
rect 1366 1458 1370 1462
rect 1326 1418 1330 1422
rect 1382 1438 1386 1442
rect 1422 1488 1426 1492
rect 1358 1418 1362 1422
rect 1326 1348 1330 1352
rect 1358 1358 1362 1362
rect 1414 1448 1418 1452
rect 1406 1418 1410 1422
rect 1414 1418 1418 1422
rect 1374 1348 1378 1352
rect 1382 1348 1386 1352
rect 1342 1338 1346 1342
rect 1350 1338 1354 1342
rect 1358 1328 1362 1332
rect 1350 1318 1354 1322
rect 1334 1288 1338 1292
rect 1246 1268 1250 1272
rect 1246 1248 1250 1252
rect 1334 1268 1338 1272
rect 1342 1268 1346 1272
rect 1286 1258 1290 1262
rect 1278 1248 1282 1252
rect 1262 1228 1266 1232
rect 1238 1198 1242 1202
rect 1294 1238 1298 1242
rect 1310 1248 1314 1252
rect 1262 1188 1266 1192
rect 1238 1178 1242 1182
rect 1294 1218 1298 1222
rect 1310 1218 1314 1222
rect 1342 1248 1346 1252
rect 1350 1248 1354 1252
rect 1334 1238 1338 1242
rect 1326 1218 1330 1222
rect 1334 1218 1338 1222
rect 1310 1198 1314 1202
rect 1318 1198 1322 1202
rect 1326 1188 1330 1192
rect 1246 1158 1250 1162
rect 1262 1158 1266 1162
rect 1286 1158 1290 1162
rect 1230 1148 1234 1152
rect 1246 1148 1250 1152
rect 1238 1128 1242 1132
rect 1246 1068 1250 1072
rect 1286 1148 1290 1152
rect 1294 1138 1298 1142
rect 1302 1138 1306 1142
rect 1278 1128 1282 1132
rect 1382 1328 1386 1332
rect 1390 1298 1394 1302
rect 1374 1288 1378 1292
rect 1358 1218 1362 1222
rect 1350 1188 1354 1192
rect 1390 1228 1394 1232
rect 1390 1208 1394 1212
rect 1390 1198 1394 1202
rect 1366 1168 1370 1172
rect 1430 1448 1434 1452
rect 1430 1378 1434 1382
rect 1470 1588 1474 1592
rect 1446 1568 1450 1572
rect 1462 1558 1466 1562
rect 1446 1548 1450 1552
rect 1454 1528 1458 1532
rect 1534 1648 1538 1652
rect 1558 1648 1562 1652
rect 1518 1628 1522 1632
rect 1534 1628 1538 1632
rect 1514 1603 1518 1607
rect 1521 1603 1525 1607
rect 1494 1598 1498 1602
rect 1486 1578 1490 1582
rect 1478 1568 1482 1572
rect 1502 1558 1506 1562
rect 1518 1558 1522 1562
rect 1494 1548 1498 1552
rect 1478 1538 1482 1542
rect 1486 1538 1490 1542
rect 1526 1538 1530 1542
rect 1478 1518 1482 1522
rect 1494 1508 1498 1512
rect 1454 1468 1458 1472
rect 1470 1458 1474 1462
rect 1502 1468 1506 1472
rect 1462 1448 1466 1452
rect 1478 1448 1482 1452
rect 1598 1658 1602 1662
rect 1614 1658 1618 1662
rect 1582 1608 1586 1612
rect 1566 1578 1570 1582
rect 1558 1558 1562 1562
rect 1574 1558 1578 1562
rect 1582 1548 1586 1552
rect 1542 1528 1546 1532
rect 1550 1518 1554 1522
rect 1582 1518 1586 1522
rect 1566 1508 1570 1512
rect 1574 1508 1578 1512
rect 1542 1468 1546 1472
rect 1574 1478 1578 1482
rect 1614 1648 1618 1652
rect 1678 1728 1682 1732
rect 1646 1718 1650 1722
rect 1670 1718 1674 1722
rect 1662 1688 1666 1692
rect 1678 1688 1682 1692
rect 1638 1678 1642 1682
rect 1710 1778 1714 1782
rect 1766 1848 1770 1852
rect 1742 1798 1746 1802
rect 1734 1778 1738 1782
rect 1726 1738 1730 1742
rect 1702 1728 1706 1732
rect 1790 1808 1794 1812
rect 1798 1798 1802 1802
rect 1774 1768 1778 1772
rect 1774 1758 1778 1762
rect 1750 1738 1754 1742
rect 1750 1728 1754 1732
rect 1742 1718 1746 1722
rect 1814 1858 1818 1862
rect 1814 1848 1818 1852
rect 1814 1828 1818 1832
rect 1814 1808 1818 1812
rect 1862 1888 1866 1892
rect 2030 1948 2034 1952
rect 2038 1928 2042 1932
rect 2030 1918 2034 1922
rect 2070 2118 2074 2122
rect 2062 2108 2066 2112
rect 2054 2068 2058 2072
rect 2054 2048 2058 2052
rect 2070 2038 2074 2042
rect 2086 2158 2090 2162
rect 2102 2158 2106 2162
rect 2110 2118 2114 2122
rect 2134 2168 2138 2172
rect 2142 2168 2146 2172
rect 2142 2158 2146 2162
rect 2126 2138 2130 2142
rect 2150 2078 2154 2082
rect 2094 2068 2098 2072
rect 2102 2058 2106 2062
rect 2134 2058 2138 2062
rect 2118 2048 2122 2052
rect 2126 2048 2130 2052
rect 2198 2268 2202 2272
rect 2222 2328 2226 2332
rect 2222 2298 2226 2302
rect 2214 2278 2218 2282
rect 2214 2268 2218 2272
rect 2222 2268 2226 2272
rect 2294 2348 2298 2352
rect 2310 2348 2314 2352
rect 2326 2348 2330 2352
rect 2262 2338 2266 2342
rect 2262 2328 2266 2332
rect 2294 2318 2298 2322
rect 2246 2298 2250 2302
rect 2254 2298 2258 2302
rect 2510 2498 2514 2502
rect 2566 2508 2570 2512
rect 2614 2548 2618 2552
rect 2726 2858 2730 2862
rect 2742 2848 2746 2852
rect 2734 2828 2738 2832
rect 2910 2938 2914 2942
rect 2934 2938 2938 2942
rect 2862 2918 2866 2922
rect 2854 2908 2858 2912
rect 2886 2878 2890 2882
rect 2766 2858 2770 2862
rect 2790 2858 2794 2862
rect 2814 2858 2818 2862
rect 2822 2858 2826 2862
rect 2766 2848 2770 2852
rect 2790 2848 2794 2852
rect 2798 2848 2802 2852
rect 2710 2778 2714 2782
rect 2758 2778 2762 2782
rect 2742 2748 2746 2752
rect 2806 2778 2810 2782
rect 2798 2758 2802 2762
rect 2798 2738 2802 2742
rect 2814 2738 2818 2742
rect 2710 2708 2714 2712
rect 2766 2728 2770 2732
rect 2790 2728 2794 2732
rect 2742 2708 2746 2712
rect 2790 2718 2794 2722
rect 2726 2688 2730 2692
rect 2750 2688 2754 2692
rect 2766 2688 2770 2692
rect 2774 2688 2778 2692
rect 2742 2668 2746 2672
rect 2766 2668 2770 2672
rect 2782 2668 2786 2672
rect 2686 2658 2690 2662
rect 2694 2658 2698 2662
rect 2734 2658 2738 2662
rect 2710 2648 2714 2652
rect 2654 2638 2658 2642
rect 2718 2638 2722 2642
rect 2654 2608 2658 2612
rect 2694 2578 2698 2582
rect 2670 2558 2674 2562
rect 2590 2528 2594 2532
rect 2598 2528 2602 2532
rect 2542 2498 2546 2502
rect 2582 2498 2586 2502
rect 2598 2498 2602 2502
rect 2526 2488 2530 2492
rect 2574 2488 2578 2492
rect 2590 2488 2594 2492
rect 2630 2488 2634 2492
rect 2654 2538 2658 2542
rect 2686 2538 2690 2542
rect 2654 2528 2658 2532
rect 2726 2568 2730 2572
rect 2734 2548 2738 2552
rect 2710 2538 2714 2542
rect 2750 2538 2754 2542
rect 2646 2498 2650 2502
rect 2486 2468 2490 2472
rect 2510 2468 2514 2472
rect 2638 2468 2642 2472
rect 2478 2458 2482 2462
rect 2486 2458 2490 2462
rect 2518 2458 2522 2462
rect 2542 2458 2546 2462
rect 2382 2348 2386 2352
rect 2350 2338 2354 2342
rect 2358 2328 2362 2332
rect 2542 2438 2546 2442
rect 2538 2403 2542 2407
rect 2545 2403 2549 2407
rect 2574 2458 2578 2462
rect 2622 2458 2626 2462
rect 2678 2518 2682 2522
rect 2590 2448 2594 2452
rect 2598 2438 2602 2442
rect 2574 2418 2578 2422
rect 2510 2358 2514 2362
rect 2534 2358 2538 2362
rect 2398 2338 2402 2342
rect 2374 2318 2378 2322
rect 2382 2288 2386 2292
rect 2326 2278 2330 2282
rect 2270 2266 2274 2270
rect 2278 2268 2282 2272
rect 2310 2268 2314 2272
rect 2318 2268 2322 2272
rect 2286 2258 2290 2262
rect 2166 2228 2170 2232
rect 2174 2228 2178 2232
rect 2198 2198 2202 2202
rect 2206 2198 2210 2202
rect 2174 2158 2178 2162
rect 2206 2158 2210 2162
rect 2238 2248 2242 2252
rect 2254 2248 2258 2252
rect 2270 2228 2274 2232
rect 2270 2178 2274 2182
rect 2246 2158 2250 2162
rect 2246 2148 2250 2152
rect 2190 2138 2194 2142
rect 2230 2128 2234 2132
rect 2214 2108 2218 2112
rect 2222 2108 2226 2112
rect 2174 2098 2178 2102
rect 2198 2078 2202 2082
rect 2230 2098 2234 2102
rect 2238 2078 2242 2082
rect 2254 2128 2258 2132
rect 2166 2068 2170 2072
rect 2238 2068 2242 2072
rect 2246 2068 2250 2072
rect 2166 2058 2170 2062
rect 2174 2058 2178 2062
rect 2102 2038 2106 2042
rect 2142 2038 2146 2042
rect 2158 2038 2162 2042
rect 2102 2018 2106 2022
rect 2086 1968 2090 1972
rect 2078 1948 2082 1952
rect 2094 1948 2098 1952
rect 2054 1928 2058 1932
rect 2026 1903 2030 1907
rect 2033 1903 2037 1907
rect 1990 1888 1994 1892
rect 2006 1888 2010 1892
rect 2038 1888 2042 1892
rect 2046 1888 2050 1892
rect 1934 1878 1938 1882
rect 2022 1878 2026 1882
rect 1918 1868 1922 1872
rect 2006 1868 2010 1872
rect 1870 1858 1874 1862
rect 1886 1858 1890 1862
rect 1862 1848 1866 1852
rect 1878 1848 1882 1852
rect 1902 1838 1906 1842
rect 1862 1828 1866 1832
rect 1894 1828 1898 1832
rect 1862 1808 1866 1812
rect 1830 1778 1834 1782
rect 1838 1768 1842 1772
rect 1862 1758 1866 1762
rect 1910 1828 1914 1832
rect 1934 1778 1938 1782
rect 1974 1848 1978 1852
rect 1982 1848 1986 1852
rect 1998 1848 2002 1852
rect 2014 1848 2018 1852
rect 1990 1828 1994 1832
rect 1958 1798 1962 1802
rect 1974 1798 1978 1802
rect 1950 1768 1954 1772
rect 1838 1748 1842 1752
rect 1910 1748 1914 1752
rect 1918 1748 1922 1752
rect 1830 1738 1834 1742
rect 1782 1728 1786 1732
rect 1798 1728 1802 1732
rect 1806 1728 1810 1732
rect 1830 1728 1834 1732
rect 1774 1718 1778 1722
rect 1750 1708 1754 1712
rect 1646 1648 1650 1652
rect 1614 1578 1618 1582
rect 1630 1578 1634 1582
rect 1814 1718 1818 1722
rect 1782 1698 1786 1702
rect 1862 1738 1866 1742
rect 1846 1718 1850 1722
rect 1886 1728 1890 1732
rect 1894 1728 1898 1732
rect 1870 1708 1874 1712
rect 1878 1708 1882 1712
rect 1870 1698 1874 1702
rect 1702 1688 1706 1692
rect 1798 1688 1802 1692
rect 1726 1678 1730 1682
rect 1702 1668 1706 1672
rect 1742 1668 1746 1672
rect 1670 1658 1674 1662
rect 1702 1648 1706 1652
rect 1726 1648 1730 1652
rect 1710 1638 1714 1642
rect 1718 1618 1722 1622
rect 1678 1608 1682 1612
rect 1670 1598 1674 1602
rect 1726 1578 1730 1582
rect 1734 1578 1738 1582
rect 1662 1568 1666 1572
rect 1622 1558 1626 1562
rect 1638 1558 1642 1562
rect 1606 1548 1610 1552
rect 1550 1448 1554 1452
rect 1486 1438 1490 1442
rect 1494 1438 1498 1442
rect 1406 1318 1410 1322
rect 1438 1348 1442 1352
rect 1438 1328 1442 1332
rect 1542 1428 1546 1432
rect 1534 1408 1538 1412
rect 1514 1403 1518 1407
rect 1521 1403 1525 1407
rect 1454 1358 1458 1362
rect 1518 1358 1522 1362
rect 1422 1268 1426 1272
rect 1438 1268 1442 1272
rect 1446 1258 1450 1262
rect 1414 1248 1418 1252
rect 1422 1228 1426 1232
rect 1454 1228 1458 1232
rect 1414 1218 1418 1222
rect 1406 1188 1410 1192
rect 1414 1178 1418 1182
rect 1502 1348 1506 1352
rect 1526 1348 1530 1352
rect 1518 1318 1522 1322
rect 1510 1288 1514 1292
rect 1486 1248 1490 1252
rect 1478 1228 1482 1232
rect 1470 1208 1474 1212
rect 1462 1198 1466 1202
rect 1446 1188 1450 1192
rect 1462 1178 1466 1182
rect 1350 1138 1354 1142
rect 1366 1138 1370 1142
rect 1414 1138 1418 1142
rect 1318 1118 1322 1122
rect 1326 1118 1330 1122
rect 1286 1098 1290 1102
rect 1302 1098 1306 1102
rect 1270 1088 1274 1092
rect 1278 1088 1282 1092
rect 1206 1058 1210 1062
rect 1222 1058 1226 1062
rect 1230 1058 1234 1062
rect 1206 1048 1210 1052
rect 1198 1028 1202 1032
rect 1198 1018 1202 1022
rect 1134 988 1138 992
rect 1126 978 1130 982
rect 1110 958 1114 962
rect 1086 948 1090 952
rect 1166 968 1170 972
rect 1054 928 1058 932
rect 1046 918 1050 922
rect 1038 888 1042 892
rect 1014 858 1018 862
rect 982 808 986 812
rect 982 798 986 802
rect 958 788 962 792
rect 766 698 770 702
rect 782 698 786 702
rect 646 648 650 652
rect 702 648 706 652
rect 718 648 722 652
rect 678 638 682 642
rect 662 608 666 612
rect 654 588 658 592
rect 638 568 642 572
rect 630 558 634 562
rect 574 548 578 552
rect 478 498 482 502
rect 558 498 562 502
rect 486 488 490 492
rect 502 468 506 472
rect 550 468 554 472
rect 710 628 714 632
rect 694 618 698 622
rect 694 568 698 572
rect 694 558 698 562
rect 710 558 714 562
rect 606 538 610 542
rect 622 538 626 542
rect 654 538 658 542
rect 614 518 618 522
rect 646 518 650 522
rect 638 498 642 502
rect 622 488 626 492
rect 662 488 666 492
rect 662 478 666 482
rect 622 468 626 472
rect 542 458 546 462
rect 598 458 602 462
rect 558 448 562 452
rect 518 438 522 442
rect 526 438 530 442
rect 558 438 562 442
rect 534 428 538 432
rect 526 418 530 422
rect 482 403 486 407
rect 489 403 493 407
rect 446 378 450 382
rect 438 318 442 322
rect 582 428 586 432
rect 606 438 610 442
rect 598 398 602 402
rect 630 448 634 452
rect 686 478 690 482
rect 814 728 818 732
rect 806 668 810 672
rect 766 578 770 582
rect 790 578 794 582
rect 798 578 802 582
rect 886 738 890 742
rect 982 738 986 742
rect 870 728 874 732
rect 942 728 946 732
rect 966 728 970 732
rect 998 808 1002 812
rect 1006 758 1010 762
rect 1054 888 1058 892
rect 1094 908 1098 912
rect 1062 878 1066 882
rect 1070 878 1074 882
rect 1118 888 1122 892
rect 1102 868 1106 872
rect 1062 858 1066 862
rect 1078 858 1082 862
rect 1094 858 1098 862
rect 1118 858 1122 862
rect 1158 948 1162 952
rect 1190 988 1194 992
rect 1158 888 1162 892
rect 1166 878 1170 882
rect 1126 848 1130 852
rect 1046 838 1050 842
rect 1038 828 1042 832
rect 1046 828 1050 832
rect 1030 738 1034 742
rect 870 718 874 722
rect 878 718 882 722
rect 878 698 882 702
rect 886 698 890 702
rect 870 678 874 682
rect 830 668 834 672
rect 846 668 850 672
rect 822 608 826 612
rect 918 688 922 692
rect 926 688 930 692
rect 870 658 874 662
rect 958 708 962 712
rect 974 708 978 712
rect 958 698 962 702
rect 950 638 954 642
rect 894 628 898 632
rect 918 628 922 632
rect 966 638 970 642
rect 998 718 1002 722
rect 1038 718 1042 722
rect 1030 708 1034 712
rect 994 703 998 707
rect 1001 703 1005 707
rect 1070 798 1074 802
rect 1126 828 1130 832
rect 1118 768 1122 772
rect 1062 758 1066 762
rect 1062 738 1066 742
rect 1078 738 1082 742
rect 1126 738 1130 742
rect 1070 718 1074 722
rect 1038 688 1042 692
rect 1078 688 1082 692
rect 982 678 986 682
rect 838 588 842 592
rect 886 588 890 592
rect 902 588 906 592
rect 878 578 882 582
rect 750 568 754 572
rect 766 568 770 572
rect 806 568 810 572
rect 734 558 738 562
rect 742 548 746 552
rect 774 548 778 552
rect 726 498 730 502
rect 686 458 690 462
rect 614 408 618 412
rect 710 448 714 452
rect 710 408 714 412
rect 590 368 594 372
rect 478 358 482 362
rect 550 358 554 362
rect 454 328 458 332
rect 502 338 506 342
rect 526 338 530 342
rect 550 338 554 342
rect 574 348 578 352
rect 638 358 642 362
rect 654 358 658 362
rect 614 348 618 352
rect 654 348 658 352
rect 702 348 706 352
rect 646 338 650 342
rect 542 328 546 332
rect 566 328 570 332
rect 534 308 538 312
rect 534 298 538 302
rect 622 328 626 332
rect 574 308 578 312
rect 582 308 586 312
rect 598 308 602 312
rect 646 318 650 322
rect 462 268 466 272
rect 502 268 506 272
rect 382 168 386 172
rect 358 138 362 142
rect 374 118 378 122
rect 374 108 378 112
rect 342 88 346 92
rect 390 88 394 92
rect 414 188 418 192
rect 454 218 458 222
rect 482 203 486 207
rect 489 203 493 207
rect 446 198 450 202
rect 430 128 434 132
rect 526 248 530 252
rect 558 248 562 252
rect 622 268 626 272
rect 582 208 586 212
rect 566 198 570 202
rect 558 188 562 192
rect 462 178 466 182
rect 470 178 474 182
rect 526 178 530 182
rect 454 168 458 172
rect 438 118 442 122
rect 454 108 458 112
rect 518 158 522 162
rect 550 158 554 162
rect 614 248 618 252
rect 622 238 626 242
rect 630 238 634 242
rect 638 238 642 242
rect 590 178 594 182
rect 574 168 578 172
rect 614 208 618 212
rect 614 178 618 182
rect 630 168 634 172
rect 670 288 674 292
rect 662 278 666 282
rect 662 258 666 262
rect 750 538 754 542
rect 742 508 746 512
rect 782 488 786 492
rect 758 478 762 482
rect 766 468 770 472
rect 750 458 754 462
rect 782 458 786 462
rect 766 448 770 452
rect 734 438 738 442
rect 726 388 730 392
rect 766 378 770 382
rect 710 338 714 342
rect 694 328 698 332
rect 718 328 722 332
rect 742 328 746 332
rect 942 588 946 592
rect 910 558 914 562
rect 926 558 930 562
rect 958 558 962 562
rect 982 558 986 562
rect 846 548 850 552
rect 838 538 842 542
rect 798 528 802 532
rect 870 528 874 532
rect 806 518 810 522
rect 822 518 826 522
rect 806 508 810 512
rect 846 498 850 502
rect 870 488 874 492
rect 822 468 826 472
rect 902 548 906 552
rect 902 538 906 542
rect 894 518 898 522
rect 878 468 882 472
rect 1094 728 1098 732
rect 1150 848 1154 852
rect 1150 778 1154 782
rect 1142 768 1146 772
rect 1142 738 1146 742
rect 1150 728 1154 732
rect 1102 718 1106 722
rect 1126 718 1130 722
rect 1134 718 1138 722
rect 1006 658 1010 662
rect 1014 628 1018 632
rect 1054 638 1058 642
rect 1070 638 1074 642
rect 1118 678 1122 682
rect 1214 988 1218 992
rect 1206 948 1210 952
rect 1254 1048 1258 1052
rect 1262 1048 1266 1052
rect 1254 1028 1258 1032
rect 1278 1048 1282 1052
rect 1318 1088 1322 1092
rect 1438 1138 1442 1142
rect 1358 1128 1362 1132
rect 1366 1128 1370 1132
rect 1422 1128 1426 1132
rect 1366 1098 1370 1102
rect 1398 1098 1402 1102
rect 1374 1088 1378 1092
rect 1334 1068 1338 1072
rect 1382 1068 1386 1072
rect 1286 1038 1290 1042
rect 1262 988 1266 992
rect 1270 988 1274 992
rect 1262 968 1266 972
rect 1270 958 1274 962
rect 1318 1048 1322 1052
rect 1310 1018 1314 1022
rect 1318 1008 1322 1012
rect 1310 978 1314 982
rect 1230 948 1234 952
rect 1254 948 1258 952
rect 1206 918 1210 922
rect 1190 878 1194 882
rect 1198 868 1202 872
rect 1198 848 1202 852
rect 1198 828 1202 832
rect 1222 918 1226 922
rect 1230 908 1234 912
rect 1262 938 1266 942
rect 1278 938 1282 942
rect 1286 928 1290 932
rect 1294 928 1298 932
rect 1294 908 1298 912
rect 1246 898 1250 902
rect 1286 898 1290 902
rect 1246 888 1250 892
rect 1270 888 1274 892
rect 1278 888 1282 892
rect 1238 868 1242 872
rect 1182 808 1186 812
rect 1206 808 1210 812
rect 1174 768 1178 772
rect 1206 758 1210 762
rect 1222 828 1226 832
rect 1222 788 1226 792
rect 1254 838 1258 842
rect 1246 828 1250 832
rect 1254 828 1258 832
rect 1238 778 1242 782
rect 1246 778 1250 782
rect 1230 768 1234 772
rect 1166 738 1170 742
rect 1182 738 1186 742
rect 1206 738 1210 742
rect 1166 708 1170 712
rect 1182 708 1186 712
rect 1134 688 1138 692
rect 1158 688 1162 692
rect 1142 678 1146 682
rect 1102 638 1106 642
rect 1086 618 1090 622
rect 1038 588 1042 592
rect 1126 578 1130 582
rect 1150 578 1154 582
rect 1094 558 1098 562
rect 1110 558 1114 562
rect 1142 558 1146 562
rect 942 548 946 552
rect 1030 548 1034 552
rect 1070 548 1074 552
rect 1118 548 1122 552
rect 1126 548 1130 552
rect 926 518 930 522
rect 990 538 994 542
rect 1046 538 1050 542
rect 1086 538 1090 542
rect 1014 528 1018 532
rect 982 518 986 522
rect 966 508 970 512
rect 926 488 930 492
rect 942 488 946 492
rect 918 478 922 482
rect 958 478 962 482
rect 854 458 858 462
rect 870 458 874 462
rect 798 448 802 452
rect 782 378 786 382
rect 854 448 858 452
rect 838 438 842 442
rect 854 378 858 382
rect 886 378 890 382
rect 814 368 818 372
rect 846 358 850 362
rect 758 338 762 342
rect 774 338 778 342
rect 686 318 690 322
rect 750 318 754 322
rect 726 308 730 312
rect 774 328 778 332
rect 814 328 818 332
rect 782 308 786 312
rect 798 308 802 312
rect 838 308 842 312
rect 822 298 826 302
rect 870 368 874 372
rect 878 368 882 372
rect 942 468 946 472
rect 942 438 946 442
rect 902 368 906 372
rect 910 358 914 362
rect 934 358 938 362
rect 910 348 914 352
rect 886 338 890 342
rect 918 338 922 342
rect 934 338 938 342
rect 870 328 874 332
rect 862 308 866 312
rect 806 278 810 282
rect 846 278 850 282
rect 918 318 922 322
rect 694 268 698 272
rect 726 268 730 272
rect 742 268 746 272
rect 798 268 802 272
rect 542 148 546 152
rect 510 138 514 142
rect 574 138 578 142
rect 510 108 514 112
rect 558 108 562 112
rect 438 68 442 72
rect 478 68 482 72
rect 262 38 266 42
rect 366 48 370 52
rect 542 98 546 102
rect 638 138 642 142
rect 654 138 658 142
rect 582 128 586 132
rect 582 118 586 122
rect 550 88 554 92
rect 710 248 714 252
rect 742 248 746 252
rect 726 238 730 242
rect 758 238 762 242
rect 718 208 722 212
rect 750 208 754 212
rect 678 198 682 202
rect 790 258 794 262
rect 806 258 810 262
rect 806 248 810 252
rect 774 178 778 182
rect 758 168 762 172
rect 790 228 794 232
rect 686 158 690 162
rect 710 158 714 162
rect 726 158 730 162
rect 726 138 730 142
rect 742 138 746 142
rect 766 138 770 142
rect 670 118 674 122
rect 622 108 626 112
rect 622 98 626 102
rect 606 88 610 92
rect 542 68 546 72
rect 670 68 674 72
rect 718 128 722 132
rect 734 128 738 132
rect 902 258 906 262
rect 822 208 826 212
rect 870 238 874 242
rect 886 238 890 242
rect 846 228 850 232
rect 838 218 842 222
rect 814 178 818 182
rect 838 178 842 182
rect 814 168 818 172
rect 718 88 722 92
rect 726 88 730 92
rect 758 88 762 92
rect 686 58 690 62
rect 486 48 490 52
rect 310 38 314 42
rect 406 28 410 32
rect 438 28 442 32
rect 454 28 458 32
rect 270 8 274 12
rect 286 8 290 12
rect 482 3 486 7
rect 489 3 493 7
rect 558 48 562 52
rect 606 48 610 52
rect 606 18 610 22
rect 534 8 538 12
rect 654 48 658 52
rect 670 48 674 52
rect 806 138 810 142
rect 806 118 810 122
rect 790 108 794 112
rect 854 208 858 212
rect 822 108 826 112
rect 902 228 906 232
rect 902 208 906 212
rect 894 178 898 182
rect 870 168 874 172
rect 862 158 866 162
rect 886 158 890 162
rect 926 278 930 282
rect 942 318 946 322
rect 994 503 998 507
rect 1001 503 1005 507
rect 1014 488 1018 492
rect 982 478 986 482
rect 1094 508 1098 512
rect 1150 538 1154 542
rect 1054 488 1058 492
rect 1086 488 1090 492
rect 1102 488 1106 492
rect 1030 478 1034 482
rect 1038 478 1042 482
rect 1078 468 1082 472
rect 1062 458 1066 462
rect 990 448 994 452
rect 1030 448 1034 452
rect 1046 438 1050 442
rect 1014 368 1018 372
rect 998 348 1002 352
rect 982 338 986 342
rect 966 328 970 332
rect 998 328 1002 332
rect 994 303 998 307
rect 1001 303 1005 307
rect 958 288 962 292
rect 1062 388 1066 392
rect 1190 698 1194 702
rect 1270 758 1274 762
rect 1302 898 1306 902
rect 1342 1038 1346 1042
rect 1358 1038 1362 1042
rect 1334 998 1338 1002
rect 1318 938 1322 942
rect 1318 908 1322 912
rect 1382 1018 1386 1022
rect 1390 1018 1394 1022
rect 1366 988 1370 992
rect 1446 1098 1450 1102
rect 1430 1068 1434 1072
rect 1558 1438 1562 1442
rect 1582 1458 1586 1462
rect 1590 1458 1594 1462
rect 1558 1378 1562 1382
rect 1574 1378 1578 1382
rect 1590 1418 1594 1422
rect 1614 1538 1618 1542
rect 1630 1528 1634 1532
rect 1614 1518 1618 1522
rect 1638 1518 1642 1522
rect 1638 1488 1642 1492
rect 1646 1488 1650 1492
rect 1614 1468 1618 1472
rect 1606 1448 1610 1452
rect 1630 1448 1634 1452
rect 1646 1448 1650 1452
rect 1702 1558 1706 1562
rect 1734 1558 1738 1562
rect 1718 1548 1722 1552
rect 1678 1538 1682 1542
rect 1694 1538 1698 1542
rect 1686 1528 1690 1532
rect 1670 1508 1674 1512
rect 1686 1508 1690 1512
rect 1662 1498 1666 1502
rect 1694 1488 1698 1492
rect 1710 1488 1714 1492
rect 1678 1478 1682 1482
rect 1702 1478 1706 1482
rect 1710 1468 1714 1472
rect 1670 1448 1674 1452
rect 1702 1448 1706 1452
rect 1710 1448 1714 1452
rect 1614 1438 1618 1442
rect 1678 1438 1682 1442
rect 1694 1438 1698 1442
rect 1646 1398 1650 1402
rect 1686 1388 1690 1392
rect 1646 1378 1650 1382
rect 1670 1368 1674 1372
rect 1598 1358 1602 1362
rect 1574 1348 1578 1352
rect 1646 1348 1650 1352
rect 1574 1328 1578 1332
rect 1566 1288 1570 1292
rect 1574 1288 1578 1292
rect 1606 1318 1610 1322
rect 1590 1298 1594 1302
rect 1590 1288 1594 1292
rect 1550 1268 1554 1272
rect 1614 1288 1618 1292
rect 1566 1258 1570 1262
rect 1598 1258 1602 1262
rect 1606 1258 1610 1262
rect 1542 1248 1546 1252
rect 1574 1248 1578 1252
rect 1582 1248 1586 1252
rect 1494 1208 1498 1212
rect 1478 1168 1482 1172
rect 1486 1168 1490 1172
rect 1478 1148 1482 1152
rect 1486 1138 1490 1142
rect 1478 1128 1482 1132
rect 1470 1098 1474 1102
rect 1446 1058 1450 1062
rect 1430 1028 1434 1032
rect 1406 988 1410 992
rect 1414 968 1418 972
rect 1462 1018 1466 1022
rect 1438 998 1442 1002
rect 1446 988 1450 992
rect 1398 948 1402 952
rect 1470 948 1474 952
rect 1350 938 1354 942
rect 1334 928 1338 932
rect 1414 938 1418 942
rect 1470 938 1474 942
rect 1390 928 1394 932
rect 1398 928 1402 932
rect 1446 928 1450 932
rect 1514 1203 1518 1207
rect 1521 1203 1525 1207
rect 1534 1168 1538 1172
rect 1510 1148 1514 1152
rect 1526 1148 1530 1152
rect 1558 1208 1562 1212
rect 1566 1188 1570 1192
rect 1558 1138 1562 1142
rect 1550 1128 1554 1132
rect 1542 1088 1546 1092
rect 1550 1088 1554 1092
rect 1606 1238 1610 1242
rect 1598 1168 1602 1172
rect 1630 1328 1634 1332
rect 1654 1318 1658 1322
rect 1638 1268 1642 1272
rect 1638 1248 1642 1252
rect 1646 1248 1650 1252
rect 1694 1348 1698 1352
rect 1710 1398 1714 1402
rect 1710 1358 1714 1362
rect 1678 1328 1682 1332
rect 1686 1328 1690 1332
rect 1726 1498 1730 1502
rect 1726 1478 1730 1482
rect 1726 1468 1730 1472
rect 1822 1678 1826 1682
rect 1830 1668 1834 1672
rect 1966 1768 1970 1772
rect 1934 1728 1938 1732
rect 1918 1718 1922 1722
rect 1926 1718 1930 1722
rect 1902 1678 1906 1682
rect 1854 1668 1858 1672
rect 1870 1668 1874 1672
rect 1894 1668 1898 1672
rect 1750 1658 1754 1662
rect 1750 1608 1754 1612
rect 1822 1648 1826 1652
rect 1814 1618 1818 1622
rect 1774 1608 1778 1612
rect 1822 1608 1826 1612
rect 1758 1558 1762 1562
rect 1798 1558 1802 1562
rect 1766 1548 1770 1552
rect 1878 1618 1882 1622
rect 1958 1708 1962 1712
rect 1974 1688 1978 1692
rect 1942 1668 1946 1672
rect 1910 1658 1914 1662
rect 1934 1658 1938 1662
rect 1966 1658 1970 1662
rect 1942 1648 1946 1652
rect 1958 1648 1962 1652
rect 1910 1618 1914 1622
rect 1918 1618 1922 1622
rect 1846 1608 1850 1612
rect 1894 1608 1898 1612
rect 1838 1558 1842 1562
rect 1886 1558 1890 1562
rect 1894 1558 1898 1562
rect 1838 1548 1842 1552
rect 1774 1528 1778 1532
rect 1758 1518 1762 1522
rect 1766 1518 1770 1522
rect 1790 1518 1794 1522
rect 1758 1508 1762 1512
rect 1790 1508 1794 1512
rect 1830 1508 1834 1512
rect 1862 1528 1866 1532
rect 1862 1518 1866 1522
rect 1846 1508 1850 1512
rect 1854 1508 1858 1512
rect 1822 1498 1826 1502
rect 1774 1488 1778 1492
rect 1782 1488 1786 1492
rect 1798 1488 1802 1492
rect 1806 1488 1810 1492
rect 1742 1478 1746 1482
rect 1782 1478 1786 1482
rect 1758 1468 1762 1472
rect 1742 1458 1746 1462
rect 1726 1448 1730 1452
rect 1734 1448 1738 1452
rect 1734 1418 1738 1422
rect 1750 1398 1754 1402
rect 1726 1358 1730 1362
rect 1766 1458 1770 1462
rect 1822 1458 1826 1462
rect 1830 1458 1834 1462
rect 1782 1428 1786 1432
rect 1782 1398 1786 1402
rect 1766 1368 1770 1372
rect 1734 1348 1738 1352
rect 1758 1348 1762 1352
rect 1774 1348 1778 1352
rect 1782 1348 1786 1352
rect 1718 1338 1722 1342
rect 1766 1338 1770 1342
rect 1726 1328 1730 1332
rect 1662 1268 1666 1272
rect 1678 1268 1682 1272
rect 1710 1268 1714 1272
rect 1734 1268 1738 1272
rect 1670 1258 1674 1262
rect 1702 1258 1706 1262
rect 1774 1308 1778 1312
rect 1766 1288 1770 1292
rect 1750 1258 1754 1262
rect 1758 1258 1762 1262
rect 1630 1208 1634 1212
rect 1638 1208 1642 1212
rect 1630 1188 1634 1192
rect 1654 1188 1658 1192
rect 1670 1188 1674 1192
rect 1622 1158 1626 1162
rect 1646 1158 1650 1162
rect 1606 1148 1610 1152
rect 1630 1148 1634 1152
rect 1646 1148 1650 1152
rect 1582 1138 1586 1142
rect 1590 1138 1594 1142
rect 1638 1138 1642 1142
rect 1574 1128 1578 1132
rect 1542 1068 1546 1072
rect 1574 1068 1578 1072
rect 1510 1058 1514 1062
rect 1494 1018 1498 1022
rect 1566 1028 1570 1032
rect 1558 1018 1562 1022
rect 1502 1008 1506 1012
rect 1514 1003 1518 1007
rect 1521 1003 1525 1007
rect 1558 998 1562 1002
rect 1534 988 1538 992
rect 1518 948 1522 952
rect 1462 928 1466 932
rect 1478 928 1482 932
rect 1358 918 1362 922
rect 1454 918 1458 922
rect 1494 918 1498 922
rect 1358 908 1362 912
rect 1366 908 1370 912
rect 1350 878 1354 882
rect 1366 878 1370 882
rect 1326 868 1330 872
rect 1342 868 1346 872
rect 1310 858 1314 862
rect 1326 858 1330 862
rect 1334 858 1338 862
rect 1294 808 1298 812
rect 1406 908 1410 912
rect 1414 908 1418 912
rect 1462 908 1466 912
rect 1398 898 1402 902
rect 1382 858 1386 862
rect 1382 848 1386 852
rect 1358 838 1362 842
rect 1342 808 1346 812
rect 1406 848 1410 852
rect 1430 868 1434 872
rect 1486 898 1490 902
rect 1478 888 1482 892
rect 1518 908 1522 912
rect 1542 958 1546 962
rect 1614 1128 1618 1132
rect 1638 1128 1642 1132
rect 1590 1048 1594 1052
rect 1622 1068 1626 1072
rect 1630 1068 1634 1072
rect 1606 1058 1610 1062
rect 1582 988 1586 992
rect 1614 998 1618 1002
rect 1582 968 1586 972
rect 1606 968 1610 972
rect 1606 948 1610 952
rect 1630 1048 1634 1052
rect 1662 1118 1666 1122
rect 1662 1098 1666 1102
rect 1654 1088 1658 1092
rect 1654 1078 1658 1082
rect 1694 1228 1698 1232
rect 1798 1428 1802 1432
rect 1806 1418 1810 1422
rect 1838 1418 1842 1422
rect 1814 1388 1818 1392
rect 1822 1368 1826 1372
rect 2190 2048 2194 2052
rect 2214 2048 2218 2052
rect 2310 2248 2314 2252
rect 2382 2268 2386 2272
rect 2414 2308 2418 2312
rect 2470 2328 2474 2332
rect 2494 2328 2498 2332
rect 2502 2328 2506 2332
rect 2614 2368 2618 2372
rect 2598 2358 2602 2362
rect 2606 2358 2610 2362
rect 2590 2348 2594 2352
rect 2750 2528 2754 2532
rect 2726 2518 2730 2522
rect 2710 2508 2714 2512
rect 2694 2498 2698 2502
rect 2670 2448 2674 2452
rect 2630 2358 2634 2362
rect 2654 2358 2658 2362
rect 2566 2328 2570 2332
rect 2486 2318 2490 2322
rect 2550 2318 2554 2322
rect 2566 2318 2570 2322
rect 2454 2298 2458 2302
rect 2406 2278 2410 2282
rect 2422 2278 2426 2282
rect 2454 2278 2458 2282
rect 2430 2268 2434 2272
rect 2390 2258 2394 2262
rect 2438 2258 2442 2262
rect 2366 2248 2370 2252
rect 2422 2248 2426 2252
rect 2446 2248 2450 2252
rect 2342 2238 2346 2242
rect 2334 2208 2338 2212
rect 2430 2198 2434 2202
rect 2406 2168 2410 2172
rect 2422 2168 2426 2172
rect 2302 2158 2306 2162
rect 2342 2158 2346 2162
rect 2374 2158 2378 2162
rect 2414 2158 2418 2162
rect 2326 2148 2330 2152
rect 2278 2138 2282 2142
rect 2302 2138 2306 2142
rect 2654 2348 2658 2352
rect 2654 2338 2658 2342
rect 2702 2438 2706 2442
rect 2734 2498 2738 2502
rect 2718 2458 2722 2462
rect 2726 2448 2730 2452
rect 2758 2458 2762 2462
rect 2766 2448 2770 2452
rect 2742 2438 2746 2442
rect 2806 2688 2810 2692
rect 2878 2858 2882 2862
rect 2846 2838 2850 2842
rect 2886 2758 2890 2762
rect 2830 2738 2834 2742
rect 2846 2738 2850 2742
rect 2862 2738 2866 2742
rect 2822 2728 2826 2732
rect 2846 2708 2850 2712
rect 2830 2698 2834 2702
rect 2838 2688 2842 2692
rect 2846 2688 2850 2692
rect 2894 2738 2898 2742
rect 2870 2698 2874 2702
rect 2894 2698 2898 2702
rect 2878 2688 2882 2692
rect 2854 2678 2858 2682
rect 2870 2678 2874 2682
rect 2798 2668 2802 2672
rect 2814 2668 2818 2672
rect 2830 2668 2834 2672
rect 2942 2928 2946 2932
rect 2926 2888 2930 2892
rect 3006 3138 3010 3142
rect 2990 3118 2994 3122
rect 3038 3138 3042 3142
rect 3022 3128 3026 3132
rect 3078 3128 3082 3132
rect 3030 3118 3034 3122
rect 3094 3118 3098 3122
rect 2990 3078 2994 3082
rect 3042 3103 3046 3107
rect 3049 3103 3053 3107
rect 2990 3058 2994 3062
rect 3046 3058 3050 3062
rect 3062 3058 3066 3062
rect 3070 3058 3074 3062
rect 3070 3048 3074 3052
rect 3006 3038 3010 3042
rect 3054 3028 3058 3032
rect 2982 2998 2986 3002
rect 2982 2978 2986 2982
rect 3022 2978 3026 2982
rect 2966 2968 2970 2972
rect 2982 2958 2986 2962
rect 3014 2958 3018 2962
rect 3014 2948 3018 2952
rect 2926 2838 2930 2842
rect 2926 2768 2930 2772
rect 2910 2678 2914 2682
rect 2846 2668 2850 2672
rect 2870 2668 2874 2672
rect 2838 2658 2842 2662
rect 2862 2658 2866 2662
rect 2806 2638 2810 2642
rect 2806 2618 2810 2622
rect 2846 2648 2850 2652
rect 2902 2658 2906 2662
rect 2854 2628 2858 2632
rect 2894 2608 2898 2612
rect 2926 2728 2930 2732
rect 2966 2818 2970 2822
rect 3046 2948 3050 2952
rect 3086 3088 3090 3092
rect 3078 2978 3082 2982
rect 3118 3278 3122 3282
rect 3126 3278 3130 3282
rect 3390 3278 3394 3282
rect 3110 3268 3114 3272
rect 3318 3268 3322 3272
rect 3374 3268 3378 3272
rect 3478 3268 3482 3272
rect 3118 3258 3122 3262
rect 3182 3258 3186 3262
rect 3390 3258 3394 3262
rect 3438 3258 3442 3262
rect 3462 3258 3466 3262
rect 3118 3238 3122 3242
rect 3142 3238 3146 3242
rect 3110 3178 3114 3182
rect 3142 3158 3146 3162
rect 3198 3178 3202 3182
rect 3222 3168 3226 3172
rect 3230 3168 3234 3172
rect 3214 3158 3218 3162
rect 3174 3138 3178 3142
rect 3294 3238 3298 3242
rect 3366 3248 3370 3252
rect 3398 3248 3402 3252
rect 3454 3248 3458 3252
rect 3494 3248 3498 3252
rect 3518 3278 3522 3282
rect 3510 3268 3514 3272
rect 3518 3258 3522 3262
rect 3358 3238 3362 3242
rect 3374 3238 3378 3242
rect 3398 3238 3402 3242
rect 3350 3168 3354 3172
rect 3270 3158 3274 3162
rect 3302 3158 3306 3162
rect 3334 3158 3338 3162
rect 3246 3148 3250 3152
rect 3182 3108 3186 3112
rect 3238 3108 3242 3112
rect 3174 3088 3178 3092
rect 3214 3088 3218 3092
rect 3326 3128 3330 3132
rect 3358 3158 3362 3162
rect 3358 3138 3362 3142
rect 3382 3158 3386 3162
rect 3414 3138 3418 3142
rect 3382 3128 3386 3132
rect 3398 3128 3402 3132
rect 3350 3118 3354 3122
rect 3382 3118 3386 3122
rect 3318 3088 3322 3092
rect 3334 3088 3338 3092
rect 3470 3228 3474 3232
rect 3430 3188 3434 3192
rect 3422 3108 3426 3112
rect 3342 3078 3346 3082
rect 3166 3068 3170 3072
rect 3254 3068 3258 3072
rect 3126 3059 3130 3063
rect 3126 3048 3130 3052
rect 3190 3048 3194 3052
rect 3214 3058 3218 3062
rect 3246 3048 3250 3052
rect 3198 3038 3202 3042
rect 3222 3038 3226 3042
rect 3318 3038 3322 3042
rect 3334 3038 3338 3042
rect 3246 2958 3250 2962
rect 3262 2958 3266 2962
rect 3278 2958 3282 2962
rect 3086 2948 3090 2952
rect 3102 2948 3106 2952
rect 3110 2948 3114 2952
rect 3158 2948 3162 2952
rect 3038 2938 3042 2942
rect 3062 2938 3066 2942
rect 3078 2938 3082 2942
rect 3102 2938 3106 2942
rect 3054 2918 3058 2922
rect 3042 2903 3046 2907
rect 3049 2903 3053 2907
rect 3014 2878 3018 2882
rect 3054 2878 3058 2882
rect 2990 2868 2994 2872
rect 3086 2888 3090 2892
rect 3078 2878 3082 2882
rect 3070 2868 3074 2872
rect 3022 2848 3026 2852
rect 2982 2818 2986 2822
rect 2974 2798 2978 2802
rect 3030 2798 3034 2802
rect 3006 2778 3010 2782
rect 3014 2768 3018 2772
rect 2982 2748 2986 2752
rect 2998 2748 3002 2752
rect 3022 2748 3026 2752
rect 2934 2708 2938 2712
rect 2950 2718 2954 2722
rect 2950 2708 2954 2712
rect 2990 2738 2994 2742
rect 2974 2708 2978 2712
rect 2982 2698 2986 2702
rect 2942 2678 2946 2682
rect 2982 2678 2986 2682
rect 3030 2728 3034 2732
rect 3022 2708 3026 2712
rect 2998 2668 3002 2672
rect 3014 2668 3018 2672
rect 2918 2598 2922 2602
rect 2854 2588 2858 2592
rect 2886 2588 2890 2592
rect 2814 2578 2818 2582
rect 2966 2618 2970 2622
rect 2942 2608 2946 2612
rect 2966 2608 2970 2612
rect 2934 2598 2938 2602
rect 2926 2578 2930 2582
rect 2894 2568 2898 2572
rect 2814 2558 2818 2562
rect 2918 2558 2922 2562
rect 2878 2548 2882 2552
rect 2814 2538 2818 2542
rect 2838 2538 2842 2542
rect 2838 2518 2842 2522
rect 2814 2468 2818 2472
rect 2782 2448 2786 2452
rect 2806 2448 2810 2452
rect 2814 2448 2818 2452
rect 2790 2438 2794 2442
rect 2774 2418 2778 2422
rect 2846 2498 2850 2502
rect 2862 2498 2866 2502
rect 2886 2488 2890 2492
rect 2958 2578 2962 2582
rect 2934 2498 2938 2502
rect 2950 2508 2954 2512
rect 2902 2468 2906 2472
rect 2894 2458 2898 2462
rect 2966 2468 2970 2472
rect 2950 2458 2954 2462
rect 2854 2448 2858 2452
rect 2918 2448 2922 2452
rect 2950 2448 2954 2452
rect 2838 2438 2842 2442
rect 2830 2398 2834 2402
rect 2718 2388 2722 2392
rect 2782 2368 2786 2372
rect 2830 2368 2834 2372
rect 2742 2358 2746 2362
rect 2822 2358 2826 2362
rect 2678 2348 2682 2352
rect 2742 2348 2746 2352
rect 2598 2328 2602 2332
rect 2646 2328 2650 2332
rect 2670 2328 2674 2332
rect 2694 2328 2698 2332
rect 2582 2298 2586 2302
rect 2590 2298 2594 2302
rect 2646 2298 2650 2302
rect 2502 2278 2506 2282
rect 2574 2278 2578 2282
rect 2494 2238 2498 2242
rect 2462 2158 2466 2162
rect 2622 2288 2626 2292
rect 2606 2278 2610 2282
rect 2574 2268 2578 2272
rect 2518 2208 2522 2212
rect 2538 2203 2542 2207
rect 2545 2203 2549 2207
rect 2518 2168 2522 2172
rect 2542 2168 2546 2172
rect 2390 2138 2394 2142
rect 2414 2138 2418 2142
rect 2502 2138 2506 2142
rect 2526 2138 2530 2142
rect 2366 2128 2370 2132
rect 2326 2118 2330 2122
rect 2422 2118 2426 2122
rect 2270 2108 2274 2112
rect 2278 2108 2282 2112
rect 2326 2108 2330 2112
rect 2294 2078 2298 2082
rect 2310 2078 2314 2082
rect 2350 2098 2354 2102
rect 2382 2078 2386 2082
rect 2390 2078 2394 2082
rect 2406 2078 2410 2082
rect 2286 2068 2290 2072
rect 2318 2068 2322 2072
rect 2438 2078 2442 2082
rect 2462 2118 2466 2122
rect 2486 2078 2490 2082
rect 2382 2058 2386 2062
rect 2398 2058 2402 2062
rect 2254 2038 2258 2042
rect 2302 2048 2306 2052
rect 2350 2048 2354 2052
rect 2366 2048 2370 2052
rect 2286 2038 2290 2042
rect 2206 1978 2210 1982
rect 2254 1978 2258 1982
rect 2110 1968 2114 1972
rect 2158 1968 2162 1972
rect 2150 1958 2154 1962
rect 2174 1958 2178 1962
rect 2118 1948 2122 1952
rect 2086 1928 2090 1932
rect 2094 1918 2098 1922
rect 2102 1918 2106 1922
rect 2062 1908 2066 1912
rect 2078 1908 2082 1912
rect 2078 1848 2082 1852
rect 2094 1838 2098 1842
rect 2078 1798 2082 1802
rect 2086 1798 2090 1802
rect 1998 1778 2002 1782
rect 2006 1768 2010 1772
rect 1990 1728 1994 1732
rect 1998 1708 2002 1712
rect 1982 1668 1986 1672
rect 2054 1758 2058 1762
rect 2062 1758 2066 1762
rect 2038 1748 2042 1752
rect 2046 1738 2050 1742
rect 2030 1728 2034 1732
rect 2026 1703 2030 1707
rect 2033 1703 2037 1707
rect 2094 1768 2098 1772
rect 2054 1698 2058 1702
rect 2062 1678 2066 1682
rect 1982 1648 1986 1652
rect 1974 1568 1978 1572
rect 2006 1568 2010 1572
rect 2022 1568 2026 1572
rect 2030 1568 2034 1572
rect 1934 1548 1938 1552
rect 1894 1528 1898 1532
rect 1870 1508 1874 1512
rect 1918 1528 1922 1532
rect 1910 1498 1914 1502
rect 1966 1548 1970 1552
rect 1942 1528 1946 1532
rect 1902 1478 1906 1482
rect 1854 1468 1858 1472
rect 1862 1468 1866 1472
rect 1854 1428 1858 1432
rect 1918 1458 1922 1462
rect 1878 1428 1882 1432
rect 1870 1408 1874 1412
rect 1918 1438 1922 1442
rect 1926 1438 1930 1442
rect 1902 1378 1906 1382
rect 1886 1368 1890 1372
rect 1918 1408 1922 1412
rect 1934 1408 1938 1412
rect 1918 1398 1922 1402
rect 1990 1528 1994 1532
rect 1990 1518 1994 1522
rect 1950 1508 1954 1512
rect 1974 1508 1978 1512
rect 1990 1508 1994 1512
rect 2022 1548 2026 1552
rect 2046 1648 2050 1652
rect 2022 1528 2026 1532
rect 2038 1528 2042 1532
rect 2026 1503 2030 1507
rect 2033 1503 2037 1507
rect 2014 1498 2018 1502
rect 2078 1728 2082 1732
rect 2078 1708 2082 1712
rect 2134 1938 2138 1942
rect 2166 1938 2170 1942
rect 2150 1928 2154 1932
rect 2118 1908 2122 1912
rect 2182 1928 2186 1932
rect 2158 1908 2162 1912
rect 2134 1898 2138 1902
rect 2190 1908 2194 1912
rect 2230 1958 2234 1962
rect 2262 1958 2266 1962
rect 2230 1938 2234 1942
rect 2214 1928 2218 1932
rect 2206 1908 2210 1912
rect 2198 1898 2202 1902
rect 2214 1898 2218 1902
rect 2206 1878 2210 1882
rect 2142 1868 2146 1872
rect 2174 1868 2178 1872
rect 2118 1858 2122 1862
rect 2142 1858 2146 1862
rect 2110 1798 2114 1802
rect 2118 1768 2122 1772
rect 2102 1758 2106 1762
rect 2118 1758 2122 1762
rect 2150 1798 2154 1802
rect 2150 1788 2154 1792
rect 2118 1748 2122 1752
rect 2142 1748 2146 1752
rect 2102 1738 2106 1742
rect 2126 1738 2130 1742
rect 2142 1738 2146 1742
rect 2158 1738 2162 1742
rect 2110 1728 2114 1732
rect 2166 1728 2170 1732
rect 2190 1788 2194 1792
rect 2238 1928 2242 1932
rect 2254 1928 2258 1932
rect 2270 1928 2274 1932
rect 2246 1908 2250 1912
rect 2294 2018 2298 2022
rect 2318 1958 2322 1962
rect 2430 2048 2434 2052
rect 2462 2048 2466 2052
rect 2486 2048 2490 2052
rect 2406 2038 2410 2042
rect 2414 2038 2418 2042
rect 2454 2038 2458 2042
rect 2478 2038 2482 2042
rect 2374 1958 2378 1962
rect 2390 1958 2394 1962
rect 2478 2028 2482 2032
rect 2414 2008 2418 2012
rect 2446 2008 2450 2012
rect 2358 1948 2362 1952
rect 2390 1948 2394 1952
rect 2318 1938 2322 1942
rect 2334 1938 2338 1942
rect 2294 1928 2298 1932
rect 2238 1888 2242 1892
rect 2246 1888 2250 1892
rect 2294 1888 2298 1892
rect 2326 1928 2330 1932
rect 2326 1888 2330 1892
rect 2238 1868 2242 1872
rect 2278 1858 2282 1862
rect 2294 1858 2298 1862
rect 2270 1848 2274 1852
rect 2262 1828 2266 1832
rect 2254 1788 2258 1792
rect 2222 1778 2226 1782
rect 2206 1758 2210 1762
rect 2198 1748 2202 1752
rect 2182 1738 2186 1742
rect 2174 1718 2178 1722
rect 2198 1718 2202 1722
rect 2126 1708 2130 1712
rect 2166 1708 2170 1712
rect 2174 1708 2178 1712
rect 2094 1698 2098 1702
rect 2118 1698 2122 1702
rect 2134 1698 2138 1702
rect 2198 1698 2202 1702
rect 2126 1688 2130 1692
rect 2150 1688 2154 1692
rect 2166 1688 2170 1692
rect 2078 1678 2082 1682
rect 2078 1648 2082 1652
rect 2054 1558 2058 1562
rect 2094 1548 2098 1552
rect 2086 1528 2090 1532
rect 2110 1648 2114 1652
rect 2118 1648 2122 1652
rect 2230 1758 2234 1762
rect 2214 1748 2218 1752
rect 2254 1738 2258 1742
rect 2214 1678 2218 1682
rect 2230 1678 2234 1682
rect 2182 1668 2186 1672
rect 2270 1788 2274 1792
rect 2278 1748 2282 1752
rect 2270 1738 2274 1742
rect 2302 1848 2306 1852
rect 2310 1808 2314 1812
rect 2334 1878 2338 1882
rect 2350 1878 2354 1882
rect 2342 1868 2346 1872
rect 2326 1848 2330 1852
rect 2374 1918 2378 1922
rect 2366 1858 2370 1862
rect 2342 1828 2346 1832
rect 2334 1808 2338 1812
rect 2334 1788 2338 1792
rect 2318 1748 2322 1752
rect 2302 1738 2306 1742
rect 2278 1698 2282 1702
rect 2310 1728 2314 1732
rect 2366 1778 2370 1782
rect 2342 1708 2346 1712
rect 2358 1728 2362 1732
rect 2366 1698 2370 1702
rect 2350 1688 2354 1692
rect 2270 1678 2274 1682
rect 2406 1888 2410 1892
rect 2422 1998 2426 2002
rect 2462 1988 2466 1992
rect 2462 1978 2466 1982
rect 2510 2098 2514 2102
rect 2534 2098 2538 2102
rect 2566 2198 2570 2202
rect 2502 2078 2506 2082
rect 2518 2078 2522 2082
rect 2558 2078 2562 2082
rect 2502 2018 2506 2022
rect 2494 2008 2498 2012
rect 2486 1958 2490 1962
rect 2454 1908 2458 1912
rect 2494 1908 2498 1912
rect 2494 1898 2498 1902
rect 2534 2018 2538 2022
rect 2518 2008 2522 2012
rect 2558 2008 2562 2012
rect 2538 2003 2542 2007
rect 2545 2003 2549 2007
rect 2518 1998 2522 2002
rect 2606 2248 2610 2252
rect 2598 2158 2602 2162
rect 2638 2268 2642 2272
rect 2638 2238 2642 2242
rect 2678 2298 2682 2302
rect 2750 2328 2754 2332
rect 2726 2308 2730 2312
rect 2686 2288 2690 2292
rect 2710 2288 2714 2292
rect 2662 2278 2666 2282
rect 2702 2278 2706 2282
rect 2734 2278 2738 2282
rect 2742 2268 2746 2272
rect 2678 2258 2682 2262
rect 2702 2258 2706 2262
rect 2718 2258 2722 2262
rect 2654 2168 2658 2172
rect 2606 2148 2610 2152
rect 2654 2148 2658 2152
rect 2582 2118 2586 2122
rect 2590 2048 2594 2052
rect 2606 2098 2610 2102
rect 2606 2088 2610 2092
rect 2606 2068 2610 2072
rect 2630 2138 2634 2142
rect 2806 2328 2810 2332
rect 2782 2298 2786 2302
rect 2838 2328 2842 2332
rect 2822 2308 2826 2312
rect 2758 2278 2762 2282
rect 2766 2278 2770 2282
rect 2806 2278 2810 2282
rect 2814 2278 2818 2282
rect 2758 2268 2762 2272
rect 2750 2258 2754 2262
rect 2766 2258 2770 2262
rect 2702 2248 2706 2252
rect 2734 2248 2738 2252
rect 2766 2248 2770 2252
rect 2742 2238 2746 2242
rect 2758 2218 2762 2222
rect 2718 2178 2722 2182
rect 2686 2148 2690 2152
rect 2750 2148 2754 2152
rect 2774 2208 2778 2212
rect 2798 2208 2802 2212
rect 2870 2438 2874 2442
rect 2894 2418 2898 2422
rect 2870 2368 2874 2372
rect 2966 2438 2970 2442
rect 2982 2658 2986 2662
rect 3070 2758 3074 2762
rect 3086 2848 3090 2852
rect 3102 2868 3106 2872
rect 3134 2938 3138 2942
rect 3150 2938 3154 2942
rect 3142 2928 3146 2932
rect 3174 2928 3178 2932
rect 3126 2918 3130 2922
rect 3158 2918 3162 2922
rect 3118 2888 3122 2892
rect 3118 2878 3122 2882
rect 3126 2868 3130 2872
rect 3094 2838 3098 2842
rect 3110 2838 3114 2842
rect 3086 2788 3090 2792
rect 3086 2738 3090 2742
rect 3054 2728 3058 2732
rect 3038 2718 3042 2722
rect 3042 2703 3046 2707
rect 3049 2703 3053 2707
rect 3038 2688 3042 2692
rect 3110 2768 3114 2772
rect 3118 2738 3122 2742
rect 3102 2698 3106 2702
rect 3078 2668 3082 2672
rect 2982 2648 2986 2652
rect 2998 2648 3002 2652
rect 3006 2588 3010 2592
rect 3038 2588 3042 2592
rect 3014 2568 3018 2572
rect 3006 2548 3010 2552
rect 3046 2568 3050 2572
rect 3086 2648 3090 2652
rect 3078 2578 3082 2582
rect 3070 2558 3074 2562
rect 3022 2528 3026 2532
rect 3062 2528 3066 2532
rect 2998 2518 3002 2522
rect 3014 2508 3018 2512
rect 2998 2478 3002 2482
rect 3042 2503 3046 2507
rect 3049 2503 3053 2507
rect 3030 2488 3034 2492
rect 2990 2468 2994 2472
rect 3038 2468 3042 2472
rect 3030 2458 3034 2462
rect 2982 2448 2986 2452
rect 3070 2468 3074 2472
rect 3118 2638 3122 2642
rect 3110 2578 3114 2582
rect 3102 2558 3106 2562
rect 3230 2948 3234 2952
rect 3254 2948 3258 2952
rect 3302 2948 3306 2952
rect 3190 2938 3194 2942
rect 3206 2928 3210 2932
rect 3198 2918 3202 2922
rect 3294 2938 3298 2942
rect 3254 2928 3258 2932
rect 3278 2928 3282 2932
rect 3182 2908 3186 2912
rect 3214 2908 3218 2912
rect 3246 2908 3250 2912
rect 3182 2878 3186 2882
rect 3206 2878 3210 2882
rect 3270 2918 3274 2922
rect 3230 2878 3234 2882
rect 3246 2868 3250 2872
rect 3182 2858 3186 2862
rect 3198 2858 3202 2862
rect 3174 2828 3178 2832
rect 3206 2818 3210 2822
rect 3150 2808 3154 2812
rect 3158 2808 3162 2812
rect 3174 2808 3178 2812
rect 3134 2758 3138 2762
rect 3166 2758 3170 2762
rect 3142 2748 3146 2752
rect 3134 2658 3138 2662
rect 3134 2648 3138 2652
rect 3182 2758 3186 2762
rect 3190 2758 3194 2762
rect 3214 2808 3218 2812
rect 3262 2858 3266 2862
rect 3222 2768 3226 2772
rect 3238 2758 3242 2762
rect 3238 2748 3242 2752
rect 3190 2728 3194 2732
rect 3198 2728 3202 2732
rect 3158 2708 3162 2712
rect 3150 2698 3154 2702
rect 3198 2718 3202 2722
rect 3174 2698 3178 2702
rect 3206 2688 3210 2692
rect 3182 2668 3186 2672
rect 3198 2668 3202 2672
rect 3150 2658 3154 2662
rect 3150 2638 3154 2642
rect 3142 2588 3146 2592
rect 3206 2598 3210 2602
rect 3198 2578 3202 2582
rect 3198 2568 3202 2572
rect 3182 2558 3186 2562
rect 3150 2548 3154 2552
rect 3126 2538 3130 2542
rect 3150 2538 3154 2542
rect 3142 2528 3146 2532
rect 3174 2528 3178 2532
rect 3110 2518 3114 2522
rect 3142 2518 3146 2522
rect 3182 2518 3186 2522
rect 3030 2438 3034 2442
rect 3062 2438 3066 2442
rect 2974 2408 2978 2412
rect 2934 2378 2938 2382
rect 2950 2368 2954 2372
rect 2918 2358 2922 2362
rect 2966 2358 2970 2362
rect 2870 2348 2874 2352
rect 2910 2348 2914 2352
rect 2942 2348 2946 2352
rect 2950 2348 2954 2352
rect 2934 2338 2938 2342
rect 2942 2338 2946 2342
rect 2862 2328 2866 2332
rect 2886 2328 2890 2332
rect 2870 2318 2874 2322
rect 2854 2308 2858 2312
rect 2878 2308 2882 2312
rect 2918 2308 2922 2312
rect 2854 2288 2858 2292
rect 2838 2218 2842 2222
rect 2814 2198 2818 2202
rect 2806 2168 2810 2172
rect 2822 2168 2826 2172
rect 2774 2158 2778 2162
rect 2830 2158 2834 2162
rect 2782 2148 2786 2152
rect 2830 2148 2834 2152
rect 2702 2138 2706 2142
rect 2726 2138 2730 2142
rect 2630 2128 2634 2132
rect 2670 2128 2674 2132
rect 2646 2108 2650 2112
rect 2678 2078 2682 2082
rect 2678 2058 2682 2062
rect 2590 2018 2594 2022
rect 2598 2018 2602 2022
rect 2550 1938 2554 1942
rect 2606 1958 2610 1962
rect 2694 2128 2698 2132
rect 2718 2098 2722 2102
rect 2790 2128 2794 2132
rect 2750 2108 2754 2112
rect 2742 2098 2746 2102
rect 2710 2088 2714 2092
rect 2734 2078 2738 2082
rect 2798 2098 2802 2102
rect 2790 2088 2794 2092
rect 2758 2078 2762 2082
rect 2782 2078 2786 2082
rect 2766 2058 2770 2062
rect 2686 2048 2690 2052
rect 2750 2048 2754 2052
rect 2758 2048 2762 2052
rect 2814 2048 2818 2052
rect 2654 2038 2658 2042
rect 2718 2038 2722 2042
rect 2766 2038 2770 2042
rect 2806 2038 2810 2042
rect 2686 1998 2690 2002
rect 2678 1958 2682 1962
rect 2654 1948 2658 1952
rect 2566 1928 2570 1932
rect 2574 1908 2578 1912
rect 2454 1868 2458 1872
rect 2590 1878 2594 1882
rect 2526 1858 2530 1862
rect 2486 1848 2490 1852
rect 2430 1838 2434 1842
rect 2414 1808 2418 1812
rect 2414 1798 2418 1802
rect 2390 1778 2394 1782
rect 2390 1748 2394 1752
rect 2390 1708 2394 1712
rect 2382 1698 2386 1702
rect 2254 1668 2258 1672
rect 2166 1658 2170 1662
rect 2182 1648 2186 1652
rect 2142 1618 2146 1622
rect 2150 1618 2154 1622
rect 2134 1578 2138 1582
rect 2142 1578 2146 1582
rect 2286 1658 2290 1662
rect 2238 1608 2242 1612
rect 2270 1638 2274 1642
rect 2278 1628 2282 1632
rect 2254 1578 2258 1582
rect 2174 1568 2178 1572
rect 2182 1568 2186 1572
rect 2214 1568 2218 1572
rect 2230 1568 2234 1572
rect 2134 1558 2138 1562
rect 2110 1548 2114 1552
rect 2150 1548 2154 1552
rect 2110 1518 2114 1522
rect 2078 1508 2082 1512
rect 2126 1538 2130 1542
rect 2190 1548 2194 1552
rect 2190 1538 2194 1542
rect 2262 1538 2266 1542
rect 2214 1528 2218 1532
rect 2134 1508 2138 1512
rect 2102 1498 2106 1502
rect 2118 1498 2122 1502
rect 2166 1498 2170 1502
rect 2190 1488 2194 1492
rect 2206 1488 2210 1492
rect 1966 1478 1970 1482
rect 1998 1478 2002 1482
rect 1958 1438 1962 1442
rect 2046 1468 2050 1472
rect 1998 1458 2002 1462
rect 2006 1448 2010 1452
rect 1990 1438 1994 1442
rect 1958 1428 1962 1432
rect 1998 1428 2002 1432
rect 1950 1408 1954 1412
rect 1942 1368 1946 1372
rect 1950 1368 1954 1372
rect 1870 1358 1874 1362
rect 1894 1358 1898 1362
rect 1910 1358 1914 1362
rect 1942 1358 1946 1362
rect 1902 1348 1906 1352
rect 1918 1348 1922 1352
rect 1830 1328 1834 1332
rect 1846 1328 1850 1332
rect 1886 1328 1890 1332
rect 1918 1328 1922 1332
rect 1934 1328 1938 1332
rect 1806 1318 1810 1322
rect 1942 1318 1946 1322
rect 1878 1308 1882 1312
rect 1886 1308 1890 1312
rect 1894 1308 1898 1312
rect 1934 1308 1938 1312
rect 1854 1298 1858 1302
rect 1806 1288 1810 1292
rect 1798 1268 1802 1272
rect 1750 1228 1754 1232
rect 1758 1178 1762 1182
rect 1686 1158 1690 1162
rect 1718 1158 1722 1162
rect 1750 1158 1754 1162
rect 1798 1188 1802 1192
rect 1774 1158 1778 1162
rect 1694 1148 1698 1152
rect 1726 1148 1730 1152
rect 1742 1148 1746 1152
rect 1758 1148 1762 1152
rect 1702 1138 1706 1142
rect 1726 1138 1730 1142
rect 1702 1128 1706 1132
rect 1750 1138 1754 1142
rect 1750 1128 1754 1132
rect 1686 1088 1690 1092
rect 1670 1078 1674 1082
rect 1678 1068 1682 1072
rect 1694 1068 1698 1072
rect 1654 1048 1658 1052
rect 1670 1048 1674 1052
rect 1670 1008 1674 1012
rect 1718 1098 1722 1102
rect 1726 1078 1730 1082
rect 1734 1078 1738 1082
rect 1718 1068 1722 1072
rect 1702 1048 1706 1052
rect 1694 1038 1698 1042
rect 1710 1038 1714 1042
rect 1830 1278 1834 1282
rect 1846 1278 1850 1282
rect 1870 1278 1874 1282
rect 1910 1298 1914 1302
rect 1926 1288 1930 1292
rect 1838 1268 1842 1272
rect 1822 1258 1826 1262
rect 1870 1258 1874 1262
rect 1878 1258 1882 1262
rect 1902 1268 1906 1272
rect 1894 1258 1898 1262
rect 1902 1258 1906 1262
rect 1822 1248 1826 1252
rect 1966 1418 1970 1422
rect 1950 1298 1954 1302
rect 1950 1288 1954 1292
rect 1998 1408 2002 1412
rect 1974 1368 1978 1372
rect 1974 1348 1978 1352
rect 1982 1338 1986 1342
rect 1990 1328 1994 1332
rect 1990 1318 1994 1322
rect 1974 1298 1978 1302
rect 1966 1278 1970 1282
rect 1942 1268 1946 1272
rect 1950 1268 1954 1272
rect 1814 1238 1818 1242
rect 1830 1228 1834 1232
rect 2078 1458 2082 1462
rect 2102 1468 2106 1472
rect 2118 1468 2122 1472
rect 2150 1468 2154 1472
rect 2094 1448 2098 1452
rect 2086 1438 2090 1442
rect 2070 1428 2074 1432
rect 2086 1398 2090 1402
rect 2070 1388 2074 1392
rect 2014 1378 2018 1382
rect 2046 1368 2050 1372
rect 2014 1358 2018 1362
rect 2062 1348 2066 1352
rect 2038 1328 2042 1332
rect 2062 1328 2066 1332
rect 2110 1458 2114 1462
rect 2126 1458 2130 1462
rect 2118 1448 2122 1452
rect 2142 1448 2146 1452
rect 2110 1408 2114 1412
rect 2102 1378 2106 1382
rect 2102 1368 2106 1372
rect 2150 1388 2154 1392
rect 2110 1358 2114 1362
rect 2102 1348 2106 1352
rect 2174 1468 2178 1472
rect 2174 1448 2178 1452
rect 2174 1398 2178 1402
rect 2182 1388 2186 1392
rect 2214 1478 2218 1482
rect 2294 1648 2298 1652
rect 2302 1628 2306 1632
rect 2310 1628 2314 1632
rect 2342 1628 2346 1632
rect 2326 1598 2330 1602
rect 2310 1588 2314 1592
rect 2302 1558 2306 1562
rect 2310 1538 2314 1542
rect 2238 1528 2242 1532
rect 2278 1528 2282 1532
rect 2286 1528 2290 1532
rect 2230 1498 2234 1502
rect 2278 1478 2282 1482
rect 2206 1458 2210 1462
rect 2214 1458 2218 1462
rect 2246 1458 2250 1462
rect 2198 1448 2202 1452
rect 2198 1368 2202 1372
rect 2182 1358 2186 1362
rect 2118 1338 2122 1342
rect 2078 1328 2082 1332
rect 2094 1328 2098 1332
rect 2070 1318 2074 1322
rect 2026 1303 2030 1307
rect 2033 1303 2037 1307
rect 2086 1298 2090 1302
rect 2110 1328 2114 1332
rect 2126 1328 2130 1332
rect 2118 1308 2122 1312
rect 2030 1278 2034 1282
rect 2078 1278 2082 1282
rect 1998 1268 2002 1272
rect 2086 1268 2090 1272
rect 1990 1228 1994 1232
rect 1886 1218 1890 1222
rect 1966 1218 1970 1222
rect 1830 1208 1834 1212
rect 1838 1208 1842 1212
rect 1838 1198 1842 1202
rect 1846 1188 1850 1192
rect 1854 1188 1858 1192
rect 1814 1158 1818 1162
rect 1806 1148 1810 1152
rect 1774 1138 1778 1142
rect 1798 1138 1802 1142
rect 1782 1128 1786 1132
rect 1790 1128 1794 1132
rect 1830 1148 1834 1152
rect 1878 1178 1882 1182
rect 1862 1148 1866 1152
rect 1830 1128 1834 1132
rect 1774 1098 1778 1102
rect 1766 1078 1770 1082
rect 1774 1078 1778 1082
rect 1830 1118 1834 1122
rect 1814 1098 1818 1102
rect 1838 1088 1842 1092
rect 1806 1078 1810 1082
rect 1830 1078 1834 1082
rect 1846 1078 1850 1082
rect 1790 1068 1794 1072
rect 1758 1058 1762 1062
rect 1742 1048 1746 1052
rect 1758 1048 1762 1052
rect 1686 1008 1690 1012
rect 1718 1008 1722 1012
rect 1734 1008 1738 1012
rect 1742 1008 1746 1012
rect 1678 998 1682 1002
rect 1742 988 1746 992
rect 1646 958 1650 962
rect 1718 958 1722 962
rect 1750 958 1754 962
rect 1678 948 1682 952
rect 1694 948 1698 952
rect 1742 948 1746 952
rect 1598 938 1602 942
rect 1606 938 1610 942
rect 1630 938 1634 942
rect 1718 938 1722 942
rect 1574 908 1578 912
rect 1550 888 1554 892
rect 1494 878 1498 882
rect 1590 898 1594 902
rect 1534 868 1538 872
rect 1582 868 1586 872
rect 1422 848 1426 852
rect 1446 848 1450 852
rect 1478 848 1482 852
rect 1454 838 1458 842
rect 1366 808 1370 812
rect 1398 808 1402 812
rect 1406 808 1410 812
rect 1302 798 1306 802
rect 1318 798 1322 802
rect 1358 798 1362 802
rect 1462 808 1466 812
rect 1478 788 1482 792
rect 1310 778 1314 782
rect 1334 778 1338 782
rect 1430 778 1434 782
rect 1246 728 1250 732
rect 1254 728 1258 732
rect 1230 698 1234 702
rect 1206 678 1210 682
rect 1214 678 1218 682
rect 1302 738 1306 742
rect 1350 768 1354 772
rect 1390 768 1394 772
rect 1414 768 1418 772
rect 1334 738 1338 742
rect 1310 728 1314 732
rect 1326 728 1330 732
rect 1294 708 1298 712
rect 1350 738 1354 742
rect 1406 738 1410 742
rect 1422 738 1426 742
rect 1374 728 1378 732
rect 1398 698 1402 702
rect 1342 688 1346 692
rect 1238 678 1242 682
rect 1310 678 1314 682
rect 1334 678 1338 682
rect 1366 678 1370 682
rect 1390 678 1394 682
rect 1174 618 1178 622
rect 1262 668 1266 672
rect 1286 668 1290 672
rect 1222 658 1226 662
rect 1230 658 1234 662
rect 1254 658 1258 662
rect 1270 658 1274 662
rect 1294 658 1298 662
rect 1206 628 1210 632
rect 1214 628 1218 632
rect 1222 628 1226 632
rect 1286 638 1290 642
rect 1238 608 1242 612
rect 1198 578 1202 582
rect 1198 568 1202 572
rect 1294 568 1298 572
rect 1318 658 1322 662
rect 1366 658 1370 662
rect 1374 648 1378 652
rect 1342 638 1346 642
rect 1358 628 1362 632
rect 1342 608 1346 612
rect 1334 578 1338 582
rect 1318 568 1322 572
rect 1222 558 1226 562
rect 1286 558 1290 562
rect 1198 548 1202 552
rect 1246 548 1250 552
rect 1182 538 1186 542
rect 1198 528 1202 532
rect 1222 528 1226 532
rect 1206 498 1210 502
rect 1270 518 1274 522
rect 1246 508 1250 512
rect 1270 498 1274 502
rect 1158 478 1162 482
rect 1102 468 1106 472
rect 1206 468 1210 472
rect 1230 468 1234 472
rect 1318 538 1322 542
rect 1326 518 1330 522
rect 1318 508 1322 512
rect 1326 468 1330 472
rect 1094 458 1098 462
rect 1118 458 1122 462
rect 1142 458 1146 462
rect 1190 458 1194 462
rect 1286 458 1290 462
rect 1302 458 1306 462
rect 1310 458 1314 462
rect 1086 378 1090 382
rect 1030 348 1034 352
rect 1038 348 1042 352
rect 1054 348 1058 352
rect 1030 318 1034 322
rect 1022 288 1026 292
rect 1038 278 1042 282
rect 1070 358 1074 362
rect 1070 288 1074 292
rect 950 258 954 262
rect 1054 258 1058 262
rect 990 248 994 252
rect 1038 248 1042 252
rect 934 238 938 242
rect 926 218 930 222
rect 910 178 914 182
rect 862 138 866 142
rect 918 168 922 172
rect 870 108 874 112
rect 910 108 914 112
rect 862 98 866 102
rect 886 98 890 102
rect 806 68 810 72
rect 830 68 834 72
rect 766 48 770 52
rect 726 38 730 42
rect 822 58 826 62
rect 870 68 874 72
rect 926 158 930 162
rect 1046 238 1050 242
rect 998 198 1002 202
rect 1030 198 1034 202
rect 950 158 954 162
rect 950 138 954 142
rect 1046 178 1050 182
rect 1094 318 1098 322
rect 1094 288 1098 292
rect 1126 398 1130 402
rect 1158 448 1162 452
rect 1150 418 1154 422
rect 1166 418 1170 422
rect 1134 388 1138 392
rect 1110 358 1114 362
rect 1134 348 1138 352
rect 1150 348 1154 352
rect 1174 348 1178 352
rect 1174 338 1178 342
rect 1118 318 1122 322
rect 1118 298 1122 302
rect 1102 278 1106 282
rect 1110 278 1114 282
rect 1142 288 1146 292
rect 1134 278 1138 282
rect 1166 278 1170 282
rect 1254 448 1258 452
rect 1246 428 1250 432
rect 1294 428 1298 432
rect 1326 408 1330 412
rect 1198 378 1202 382
rect 1286 358 1290 362
rect 1382 578 1386 582
rect 1366 558 1370 562
rect 1494 838 1498 842
rect 1514 803 1518 807
rect 1521 803 1525 807
rect 1502 788 1506 792
rect 1526 788 1530 792
rect 1574 858 1578 862
rect 1590 848 1594 852
rect 1550 838 1554 842
rect 1566 828 1570 832
rect 1542 808 1546 812
rect 1486 768 1490 772
rect 1574 768 1578 772
rect 1446 758 1450 762
rect 1590 758 1594 762
rect 1438 708 1442 712
rect 1406 658 1410 662
rect 1470 728 1474 732
rect 1478 728 1482 732
rect 1470 678 1474 682
rect 1470 668 1474 672
rect 1550 738 1554 742
rect 1582 738 1586 742
rect 1590 738 1594 742
rect 1510 728 1514 732
rect 1542 728 1546 732
rect 1502 718 1506 722
rect 1510 678 1514 682
rect 1462 658 1466 662
rect 1494 658 1498 662
rect 1430 648 1434 652
rect 1414 598 1418 602
rect 1382 548 1386 552
rect 1342 538 1346 542
rect 1342 508 1346 512
rect 1358 508 1362 512
rect 1414 538 1418 542
rect 1438 528 1442 532
rect 1422 518 1426 522
rect 1430 498 1434 502
rect 1438 498 1442 502
rect 1406 488 1410 492
rect 1430 488 1434 492
rect 1462 648 1466 652
rect 1478 648 1482 652
rect 1486 628 1490 632
rect 1478 548 1482 552
rect 1454 538 1458 542
rect 1462 508 1466 512
rect 1478 508 1482 512
rect 1422 468 1426 472
rect 1342 458 1346 462
rect 1398 458 1402 462
rect 1414 458 1418 462
rect 1514 603 1518 607
rect 1521 603 1525 607
rect 1502 568 1506 572
rect 1518 558 1522 562
rect 1534 538 1538 542
rect 1526 528 1530 532
rect 1494 488 1498 492
rect 1510 468 1514 472
rect 1526 468 1530 472
rect 1430 448 1434 452
rect 1430 418 1434 422
rect 1446 418 1450 422
rect 1390 408 1394 412
rect 1374 398 1378 402
rect 1446 408 1450 412
rect 1398 388 1402 392
rect 1334 378 1338 382
rect 1430 368 1434 372
rect 1438 368 1442 372
rect 1406 358 1410 362
rect 1206 348 1210 352
rect 1222 348 1226 352
rect 1230 348 1234 352
rect 1254 348 1258 352
rect 1310 348 1314 352
rect 1350 348 1354 352
rect 1390 348 1394 352
rect 1182 298 1186 302
rect 1198 318 1202 322
rect 1190 288 1194 292
rect 1150 258 1154 262
rect 1182 258 1186 262
rect 1102 248 1106 252
rect 1118 248 1122 252
rect 1094 238 1098 242
rect 1126 228 1130 232
rect 1238 338 1242 342
rect 1262 338 1266 342
rect 1222 288 1226 292
rect 1278 318 1282 322
rect 1246 308 1250 312
rect 1254 308 1258 312
rect 1254 298 1258 302
rect 1246 258 1250 262
rect 1198 238 1202 242
rect 1190 228 1194 232
rect 1190 218 1194 222
rect 1134 168 1138 172
rect 1086 158 1090 162
rect 1054 138 1058 142
rect 926 128 930 132
rect 966 128 970 132
rect 982 128 986 132
rect 950 108 954 112
rect 942 98 946 102
rect 958 68 962 72
rect 846 48 850 52
rect 870 48 874 52
rect 790 38 794 42
rect 814 38 818 42
rect 702 28 706 32
rect 726 28 730 32
rect 782 28 786 32
rect 646 18 650 22
rect 662 18 666 22
rect 694 18 698 22
rect 622 8 626 12
rect 806 8 810 12
rect 886 8 890 12
rect 994 103 998 107
rect 1001 103 1005 107
rect 982 98 986 102
rect 1022 98 1026 102
rect 990 78 994 82
rect 1038 78 1042 82
rect 1054 78 1058 82
rect 1030 58 1034 62
rect 1022 48 1026 52
rect 974 8 978 12
rect 1110 138 1114 142
rect 1198 208 1202 212
rect 1230 208 1234 212
rect 1206 188 1210 192
rect 1214 168 1218 172
rect 1222 168 1226 172
rect 1158 138 1162 142
rect 1182 138 1186 142
rect 1214 138 1218 142
rect 1150 118 1154 122
rect 1174 118 1178 122
rect 1190 118 1194 122
rect 1110 108 1114 112
rect 1102 98 1106 102
rect 1070 78 1074 82
rect 1062 28 1066 32
rect 1046 8 1050 12
rect 1158 98 1162 102
rect 1126 88 1130 92
rect 1206 78 1210 82
rect 1246 148 1250 152
rect 1270 278 1274 282
rect 1286 268 1290 272
rect 1262 258 1266 262
rect 1302 258 1306 262
rect 1270 248 1274 252
rect 1286 248 1290 252
rect 1262 238 1266 242
rect 1286 228 1290 232
rect 1374 338 1378 342
rect 1382 318 1386 322
rect 1334 308 1338 312
rect 1350 308 1354 312
rect 1366 308 1370 312
rect 1326 288 1330 292
rect 1374 288 1378 292
rect 1318 278 1322 282
rect 1366 278 1370 282
rect 1342 268 1346 272
rect 1422 318 1426 322
rect 1430 308 1434 312
rect 1446 358 1450 362
rect 1486 438 1490 442
rect 1486 418 1490 422
rect 1470 388 1474 392
rect 1462 338 1466 342
rect 1326 258 1330 262
rect 1318 208 1322 212
rect 1350 178 1354 182
rect 1334 158 1338 162
rect 1342 158 1346 162
rect 1366 158 1370 162
rect 1302 148 1306 152
rect 1358 148 1362 152
rect 1262 138 1266 142
rect 1286 138 1290 142
rect 1230 128 1234 132
rect 1238 118 1242 122
rect 1262 118 1266 122
rect 1078 68 1082 72
rect 1094 68 1098 72
rect 1182 68 1186 72
rect 1238 68 1242 72
rect 1094 58 1098 62
rect 1086 38 1090 42
rect 1118 58 1122 62
rect 1214 58 1218 62
rect 1246 58 1250 62
rect 1230 48 1234 52
rect 1246 48 1250 52
rect 1342 138 1346 142
rect 1310 108 1314 112
rect 1294 78 1298 82
rect 1358 128 1362 132
rect 1350 78 1354 82
rect 1406 248 1410 252
rect 1422 258 1426 262
rect 1454 328 1458 332
rect 1470 308 1474 312
rect 1454 278 1458 282
rect 1478 278 1482 282
rect 1518 448 1522 452
rect 1514 403 1518 407
rect 1521 403 1525 407
rect 1526 348 1530 352
rect 1494 328 1498 332
rect 1526 328 1530 332
rect 1518 308 1522 312
rect 1462 268 1466 272
rect 1470 268 1474 272
rect 1486 268 1490 272
rect 1478 258 1482 262
rect 1462 248 1466 252
rect 1454 238 1458 242
rect 1446 228 1450 232
rect 1414 198 1418 202
rect 1430 198 1434 202
rect 1406 168 1410 172
rect 1446 178 1450 182
rect 1414 148 1418 152
rect 1446 148 1450 152
rect 1374 138 1378 142
rect 1390 138 1394 142
rect 1430 138 1434 142
rect 1390 128 1394 132
rect 1382 118 1386 122
rect 1398 118 1402 122
rect 1382 98 1386 102
rect 1454 128 1458 132
rect 1550 618 1554 622
rect 1550 598 1554 602
rect 1566 708 1570 712
rect 1590 678 1594 682
rect 1590 658 1594 662
rect 1574 608 1578 612
rect 1574 598 1578 602
rect 1558 578 1562 582
rect 1550 568 1554 572
rect 1614 898 1618 902
rect 1606 888 1610 892
rect 1686 928 1690 932
rect 1622 888 1626 892
rect 1654 888 1658 892
rect 1614 878 1618 882
rect 1622 878 1626 882
rect 1646 878 1650 882
rect 1614 828 1618 832
rect 1630 828 1634 832
rect 1646 828 1650 832
rect 1606 768 1610 772
rect 1670 878 1674 882
rect 1678 878 1682 882
rect 1718 918 1722 922
rect 1702 878 1706 882
rect 1662 858 1666 862
rect 1678 858 1682 862
rect 1662 848 1666 852
rect 1686 848 1690 852
rect 1734 858 1738 862
rect 1654 808 1658 812
rect 1702 808 1706 812
rect 1654 798 1658 802
rect 1638 788 1642 792
rect 1694 788 1698 792
rect 1630 768 1634 772
rect 1654 768 1658 772
rect 1662 748 1666 752
rect 1686 738 1690 742
rect 1670 728 1674 732
rect 1614 718 1618 722
rect 1654 718 1658 722
rect 1622 698 1626 702
rect 1646 698 1650 702
rect 1678 688 1682 692
rect 1718 808 1722 812
rect 1750 918 1754 922
rect 1790 1008 1794 1012
rect 1878 1128 1882 1132
rect 1862 1118 1866 1122
rect 1862 1088 1866 1092
rect 1814 1028 1818 1032
rect 1782 958 1786 962
rect 1806 958 1810 962
rect 1806 948 1810 952
rect 1790 938 1794 942
rect 1814 938 1818 942
rect 1806 908 1810 912
rect 1766 878 1770 882
rect 1798 878 1802 882
rect 1750 868 1754 872
rect 1822 868 1826 872
rect 1846 940 1850 944
rect 1958 1188 1962 1192
rect 1926 1178 1930 1182
rect 1910 1168 1914 1172
rect 1918 1168 1922 1172
rect 2022 1238 2026 1242
rect 2038 1218 2042 1222
rect 2054 1238 2058 1242
rect 2022 1208 2026 1212
rect 2046 1208 2050 1212
rect 1998 1198 2002 1202
rect 2014 1198 2018 1202
rect 1958 1158 1962 1162
rect 1966 1158 1970 1162
rect 1990 1158 1994 1162
rect 1998 1158 2002 1162
rect 1982 1148 1986 1152
rect 1990 1138 1994 1142
rect 1926 1128 1930 1132
rect 1942 1128 1946 1132
rect 1910 1118 1914 1122
rect 1934 1118 1938 1122
rect 1958 1098 1962 1102
rect 1886 1088 1890 1092
rect 1894 1088 1898 1092
rect 1878 1078 1882 1082
rect 1886 1078 1890 1082
rect 1886 1048 1890 1052
rect 1878 1038 1882 1042
rect 1878 1028 1882 1032
rect 1870 1008 1874 1012
rect 1886 968 1890 972
rect 2126 1298 2130 1302
rect 2142 1288 2146 1292
rect 2166 1328 2170 1332
rect 2134 1268 2138 1272
rect 2158 1268 2162 1272
rect 2110 1258 2114 1262
rect 2166 1248 2170 1252
rect 2102 1238 2106 1242
rect 2150 1238 2154 1242
rect 2158 1238 2162 1242
rect 2134 1228 2138 1232
rect 2150 1228 2154 1232
rect 2078 1208 2082 1212
rect 2134 1208 2138 1212
rect 2070 1198 2074 1202
rect 2046 1188 2050 1192
rect 2006 1138 2010 1142
rect 2022 1138 2026 1142
rect 1998 1128 2002 1132
rect 2006 1118 2010 1122
rect 2038 1118 2042 1122
rect 1982 1108 1986 1112
rect 2026 1103 2030 1107
rect 2033 1103 2037 1107
rect 1998 1098 2002 1102
rect 1910 1078 1914 1082
rect 1966 1078 1970 1082
rect 1974 1078 1978 1082
rect 2062 1178 2066 1182
rect 2054 1158 2058 1162
rect 2118 1188 2122 1192
rect 2126 1178 2130 1182
rect 2142 1178 2146 1182
rect 2102 1138 2106 1142
rect 2118 1138 2122 1142
rect 2070 1108 2074 1112
rect 2014 1088 2018 1092
rect 2046 1088 2050 1092
rect 1902 1068 1906 1072
rect 1902 1038 1906 1042
rect 1918 1048 1922 1052
rect 1942 1038 1946 1042
rect 1934 1008 1938 1012
rect 1902 998 1906 1002
rect 1910 998 1914 1002
rect 2062 1078 2066 1082
rect 1974 1068 1978 1072
rect 1990 1068 1994 1072
rect 2038 1068 2042 1072
rect 2046 1068 2050 1072
rect 1998 1058 2002 1062
rect 1966 1048 1970 1052
rect 1950 1018 1954 1022
rect 1982 958 1986 962
rect 1878 948 1882 952
rect 1894 948 1898 952
rect 1910 948 1914 952
rect 1974 948 1978 952
rect 1838 908 1842 912
rect 1886 908 1890 912
rect 1846 888 1850 892
rect 1926 938 1930 942
rect 1918 918 1922 922
rect 1758 858 1762 862
rect 1774 858 1778 862
rect 1830 858 1834 862
rect 1894 858 1898 862
rect 1766 838 1770 842
rect 1750 798 1754 802
rect 1838 848 1842 852
rect 1806 828 1810 832
rect 1798 788 1802 792
rect 1830 788 1834 792
rect 1814 768 1818 772
rect 1886 848 1890 852
rect 1878 798 1882 802
rect 1734 748 1738 752
rect 1830 748 1834 752
rect 1878 748 1882 752
rect 1710 738 1714 742
rect 1750 738 1754 742
rect 1718 728 1722 732
rect 1742 728 1746 732
rect 1766 728 1770 732
rect 1606 678 1610 682
rect 1662 678 1666 682
rect 1614 658 1618 662
rect 1646 658 1650 662
rect 1662 648 1666 652
rect 1598 628 1602 632
rect 1614 628 1618 632
rect 1622 618 1626 622
rect 1606 578 1610 582
rect 1598 558 1602 562
rect 1590 548 1594 552
rect 1598 538 1602 542
rect 1590 508 1594 512
rect 1550 488 1554 492
rect 1590 488 1594 492
rect 1550 418 1554 422
rect 1542 408 1546 412
rect 1542 348 1546 352
rect 1654 568 1658 572
rect 1614 508 1618 512
rect 1654 548 1658 552
rect 1638 538 1642 542
rect 1734 718 1738 722
rect 1726 688 1730 692
rect 1718 678 1722 682
rect 1694 668 1698 672
rect 1718 668 1722 672
rect 1734 668 1738 672
rect 1686 648 1690 652
rect 1750 648 1754 652
rect 1734 638 1738 642
rect 1694 628 1698 632
rect 1710 608 1714 612
rect 1750 568 1754 572
rect 1694 558 1698 562
rect 1742 558 1746 562
rect 1998 1048 2002 1052
rect 2006 998 2010 1002
rect 2086 1088 2090 1092
rect 2102 1108 2106 1112
rect 2126 1108 2130 1112
rect 2118 1088 2122 1092
rect 2094 1068 2098 1072
rect 2086 1058 2090 1062
rect 2078 1048 2082 1052
rect 2094 1048 2098 1052
rect 2070 998 2074 1002
rect 2118 1068 2122 1072
rect 2142 1138 2146 1142
rect 2110 1048 2114 1052
rect 2102 978 2106 982
rect 2046 968 2050 972
rect 2086 968 2090 972
rect 1990 948 1994 952
rect 2022 948 2026 952
rect 2054 938 2058 942
rect 2070 938 2074 942
rect 2062 928 2066 932
rect 2094 928 2098 932
rect 1934 918 1938 922
rect 1942 918 1946 922
rect 2054 918 2058 922
rect 2094 918 2098 922
rect 1950 888 1954 892
rect 1958 878 1962 882
rect 1974 878 1978 882
rect 2006 888 2010 892
rect 1934 858 1938 862
rect 1958 858 1962 862
rect 1982 858 1986 862
rect 1990 858 1994 862
rect 2046 908 2050 912
rect 2026 903 2030 907
rect 2033 903 2037 907
rect 1934 848 1938 852
rect 1966 848 1970 852
rect 1982 838 1986 842
rect 2038 838 2042 842
rect 1902 818 1906 822
rect 1934 808 1938 812
rect 1902 798 1906 802
rect 1910 798 1914 802
rect 1838 738 1842 742
rect 1862 738 1866 742
rect 1894 738 1898 742
rect 1862 718 1866 722
rect 1830 708 1834 712
rect 1790 698 1794 702
rect 1822 698 1826 702
rect 1774 688 1778 692
rect 1766 678 1770 682
rect 1774 668 1778 672
rect 1822 688 1826 692
rect 1846 688 1850 692
rect 1854 688 1858 692
rect 1886 688 1890 692
rect 1846 658 1850 662
rect 1870 638 1874 642
rect 1822 598 1826 602
rect 1910 788 1914 792
rect 1950 798 1954 802
rect 1942 788 1946 792
rect 1942 758 1946 762
rect 1998 788 2002 792
rect 2014 788 2018 792
rect 2070 868 2074 872
rect 2086 868 2090 872
rect 2070 858 2074 862
rect 2054 848 2058 852
rect 2078 848 2082 852
rect 2118 938 2122 942
rect 2158 1168 2162 1172
rect 2166 1168 2170 1172
rect 2254 1448 2258 1452
rect 2222 1388 2226 1392
rect 2230 1358 2234 1362
rect 2246 1428 2250 1432
rect 2198 1328 2202 1332
rect 2198 1308 2202 1312
rect 2206 1298 2210 1302
rect 2190 1288 2194 1292
rect 2222 1318 2226 1322
rect 2238 1318 2242 1322
rect 2222 1298 2226 1302
rect 2254 1408 2258 1412
rect 2286 1468 2290 1472
rect 2310 1488 2314 1492
rect 2294 1438 2298 1442
rect 2278 1398 2282 1402
rect 2318 1458 2322 1462
rect 2310 1398 2314 1402
rect 2358 1638 2362 1642
rect 2350 1588 2354 1592
rect 2374 1628 2378 1632
rect 2374 1558 2378 1562
rect 2358 1538 2362 1542
rect 2350 1498 2354 1502
rect 2398 1688 2402 1692
rect 2398 1678 2402 1682
rect 2414 1678 2418 1682
rect 2558 1828 2562 1832
rect 2430 1818 2434 1822
rect 2446 1818 2450 1822
rect 2494 1808 2498 1812
rect 2558 1808 2562 1812
rect 2538 1803 2542 1807
rect 2545 1803 2549 1807
rect 2454 1798 2458 1802
rect 2510 1788 2514 1792
rect 2502 1768 2506 1772
rect 2454 1758 2458 1762
rect 2438 1748 2442 1752
rect 2454 1748 2458 1752
rect 2438 1738 2442 1742
rect 2430 1728 2434 1732
rect 2462 1708 2466 1712
rect 2462 1678 2466 1682
rect 2606 1908 2610 1912
rect 2814 2018 2818 2022
rect 2742 1988 2746 1992
rect 2758 1988 2762 1992
rect 2710 1968 2714 1972
rect 2726 1958 2730 1962
rect 2638 1938 2642 1942
rect 2662 1918 2666 1922
rect 2614 1898 2618 1902
rect 2654 1888 2658 1892
rect 2694 1888 2698 1892
rect 2630 1878 2634 1882
rect 2670 1878 2674 1882
rect 2694 1878 2698 1882
rect 2622 1868 2626 1872
rect 2654 1868 2658 1872
rect 2670 1868 2674 1872
rect 2686 1868 2690 1872
rect 2662 1858 2666 1862
rect 2862 2248 2866 2252
rect 2862 2198 2866 2202
rect 2862 2148 2866 2152
rect 2838 2138 2842 2142
rect 2846 2138 2850 2142
rect 2854 2138 2858 2142
rect 2830 2098 2834 2102
rect 2846 2108 2850 2112
rect 2870 2128 2874 2132
rect 2862 2118 2866 2122
rect 2934 2298 2938 2302
rect 2926 2288 2930 2292
rect 2910 2278 2914 2282
rect 3014 2328 3018 2332
rect 2982 2298 2986 2302
rect 2998 2298 3002 2302
rect 2998 2278 3002 2282
rect 3054 2408 3058 2412
rect 3038 2348 3042 2352
rect 3054 2318 3058 2322
rect 3042 2303 3046 2307
rect 3049 2303 3053 2307
rect 3062 2268 3066 2272
rect 2902 2248 2906 2252
rect 2886 2238 2890 2242
rect 2918 2208 2922 2212
rect 2902 2188 2906 2192
rect 2934 2188 2938 2192
rect 3054 2258 3058 2262
rect 2950 2248 2954 2252
rect 2974 2218 2978 2222
rect 3038 2248 3042 2252
rect 3070 2248 3074 2252
rect 3102 2498 3106 2502
rect 3126 2498 3130 2502
rect 3118 2488 3122 2492
rect 3110 2478 3114 2482
rect 3094 2408 3098 2412
rect 3102 2398 3106 2402
rect 3094 2378 3098 2382
rect 3086 2348 3090 2352
rect 3158 2508 3162 2512
rect 3166 2488 3170 2492
rect 3198 2488 3202 2492
rect 3118 2468 3122 2472
rect 3174 2468 3178 2472
rect 3118 2458 3122 2462
rect 3142 2458 3146 2462
rect 3134 2448 3138 2452
rect 3198 2448 3202 2452
rect 3118 2428 3122 2432
rect 3182 2428 3186 2432
rect 3142 2368 3146 2372
rect 3230 2728 3234 2732
rect 3254 2778 3258 2782
rect 3262 2768 3266 2772
rect 3326 2878 3330 2882
rect 3334 2878 3338 2882
rect 3326 2868 3330 2872
rect 3350 2918 3354 2922
rect 3374 2938 3378 2942
rect 3422 2928 3426 2932
rect 3366 2908 3370 2912
rect 3398 2908 3402 2912
rect 3438 2898 3442 2902
rect 3350 2888 3354 2892
rect 3374 2888 3378 2892
rect 3446 2888 3450 2892
rect 3374 2878 3378 2882
rect 3350 2868 3354 2872
rect 3414 2868 3418 2872
rect 3438 2868 3442 2872
rect 3326 2858 3330 2862
rect 3342 2858 3346 2862
rect 3350 2858 3354 2862
rect 3294 2848 3298 2852
rect 3310 2848 3314 2852
rect 3334 2848 3338 2852
rect 3286 2838 3290 2842
rect 3318 2828 3322 2832
rect 3326 2818 3330 2822
rect 3286 2808 3290 2812
rect 3350 2838 3354 2842
rect 3406 2798 3410 2802
rect 3334 2788 3338 2792
rect 3318 2778 3322 2782
rect 3278 2758 3282 2762
rect 3286 2748 3290 2752
rect 3294 2748 3298 2752
rect 3310 2748 3314 2752
rect 3278 2728 3282 2732
rect 3246 2718 3250 2722
rect 3270 2718 3274 2722
rect 3294 2718 3298 2722
rect 3358 2758 3362 2762
rect 3342 2728 3346 2732
rect 3326 2718 3330 2722
rect 3310 2688 3314 2692
rect 3286 2678 3290 2682
rect 3270 2668 3274 2672
rect 3238 2628 3242 2632
rect 3222 2608 3226 2612
rect 3358 2738 3362 2742
rect 3446 2858 3450 2862
rect 3446 2808 3450 2812
rect 3430 2768 3434 2772
rect 3478 3198 3482 3202
rect 3502 3158 3506 3162
rect 3462 3118 3466 3122
rect 3486 2968 3490 2972
rect 3470 2948 3474 2952
rect 3486 2948 3490 2952
rect 3518 3148 3522 3152
rect 3534 3138 3538 3142
rect 3518 2978 3522 2982
rect 3518 2968 3522 2972
rect 3558 3148 3562 3152
rect 3542 2968 3546 2972
rect 3534 2948 3538 2952
rect 3542 2948 3546 2952
rect 3534 2908 3538 2912
rect 3526 2898 3530 2902
rect 3478 2878 3482 2882
rect 3494 2878 3498 2882
rect 3510 2878 3514 2882
rect 3518 2878 3522 2882
rect 3534 2878 3538 2882
rect 3478 2868 3482 2872
rect 3502 2868 3506 2872
rect 3534 2868 3538 2872
rect 3470 2858 3474 2862
rect 3494 2858 3498 2862
rect 3526 2858 3530 2862
rect 3542 2858 3546 2862
rect 3454 2798 3458 2802
rect 3510 2848 3514 2852
rect 3478 2788 3482 2792
rect 3470 2778 3474 2782
rect 3534 2778 3538 2782
rect 3478 2768 3482 2772
rect 3486 2768 3490 2772
rect 3502 2768 3506 2772
rect 3526 2758 3530 2762
rect 3542 2758 3546 2762
rect 3446 2748 3450 2752
rect 3510 2748 3514 2752
rect 3398 2738 3402 2742
rect 3406 2738 3410 2742
rect 3358 2718 3362 2722
rect 3350 2698 3354 2702
rect 3406 2708 3410 2712
rect 3366 2688 3370 2692
rect 3374 2678 3378 2682
rect 3390 2678 3394 2682
rect 3462 2738 3466 2742
rect 3478 2728 3482 2732
rect 3558 2748 3562 2752
rect 3526 2728 3530 2732
rect 3446 2718 3450 2722
rect 3518 2718 3522 2722
rect 3486 2708 3490 2712
rect 3422 2688 3426 2692
rect 3430 2688 3434 2692
rect 3478 2688 3482 2692
rect 3414 2668 3418 2672
rect 3334 2658 3338 2662
rect 3286 2648 3290 2652
rect 3286 2628 3290 2632
rect 3342 2628 3346 2632
rect 3334 2618 3338 2622
rect 3246 2578 3250 2582
rect 3342 2578 3346 2582
rect 3390 2658 3394 2662
rect 3406 2648 3410 2652
rect 3414 2648 3418 2652
rect 3374 2598 3378 2602
rect 3350 2568 3354 2572
rect 3366 2568 3370 2572
rect 3286 2548 3290 2552
rect 3318 2548 3322 2552
rect 3238 2528 3242 2532
rect 3262 2528 3266 2532
rect 3222 2468 3226 2472
rect 3254 2468 3258 2472
rect 3246 2458 3250 2462
rect 3310 2518 3314 2522
rect 3286 2508 3290 2512
rect 3310 2498 3314 2502
rect 3294 2488 3298 2492
rect 3494 2698 3498 2702
rect 3494 2678 3498 2682
rect 3558 2688 3562 2692
rect 3446 2668 3450 2672
rect 3558 2668 3562 2672
rect 3518 2638 3522 2642
rect 3406 2608 3410 2612
rect 3438 2608 3442 2612
rect 3438 2598 3442 2602
rect 3398 2568 3402 2572
rect 3422 2558 3426 2562
rect 3390 2548 3394 2552
rect 3462 2578 3466 2582
rect 3558 2578 3562 2582
rect 3374 2538 3378 2542
rect 3342 2528 3346 2532
rect 3334 2488 3338 2492
rect 3422 2518 3426 2522
rect 3374 2478 3378 2482
rect 3382 2478 3386 2482
rect 3422 2478 3426 2482
rect 3390 2468 3394 2472
rect 3414 2458 3418 2462
rect 3270 2448 3274 2452
rect 3342 2448 3346 2452
rect 3366 2448 3370 2452
rect 3390 2448 3394 2452
rect 3302 2438 3306 2442
rect 3230 2428 3234 2432
rect 3278 2428 3282 2432
rect 3246 2368 3250 2372
rect 3334 2368 3338 2372
rect 3214 2358 3218 2362
rect 3238 2358 3242 2362
rect 3254 2358 3258 2362
rect 3294 2358 3298 2362
rect 3326 2358 3330 2362
rect 3094 2338 3098 2342
rect 3126 2338 3130 2342
rect 3134 2298 3138 2302
rect 3126 2268 3130 2272
rect 3118 2258 3122 2262
rect 3094 2248 3098 2252
rect 3078 2238 3082 2242
rect 3134 2248 3138 2252
rect 3102 2218 3106 2222
rect 2998 2208 3002 2212
rect 2950 2198 2954 2202
rect 2934 2168 2938 2172
rect 2926 2158 2930 2162
rect 2942 2158 2946 2162
rect 2894 2148 2898 2152
rect 2902 2138 2906 2142
rect 2910 2128 2914 2132
rect 2918 2128 2922 2132
rect 2934 2128 2938 2132
rect 2894 2088 2898 2092
rect 2934 2088 2938 2092
rect 2886 2078 2890 2082
rect 2902 2078 2906 2082
rect 2910 2068 2914 2072
rect 2918 2068 2922 2072
rect 2918 2048 2922 2052
rect 2862 2028 2866 2032
rect 2870 2028 2874 2032
rect 2942 2038 2946 2042
rect 2974 2178 2978 2182
rect 3022 2178 3026 2182
rect 3110 2178 3114 2182
rect 2966 2158 2970 2162
rect 3006 2158 3010 2162
rect 2958 2138 2962 2142
rect 2990 2128 2994 2132
rect 2998 2128 3002 2132
rect 2966 2088 2970 2092
rect 2974 2078 2978 2082
rect 2894 2028 2898 2032
rect 2950 2028 2954 2032
rect 2878 2018 2882 2022
rect 3070 2168 3074 2172
rect 3166 2348 3170 2352
rect 3190 2348 3194 2352
rect 3166 2338 3170 2342
rect 3198 2338 3202 2342
rect 3166 2308 3170 2312
rect 3158 2278 3162 2282
rect 3158 2258 3162 2262
rect 3150 2238 3154 2242
rect 3174 2298 3178 2302
rect 3238 2338 3242 2342
rect 3230 2328 3234 2332
rect 3470 2448 3474 2452
rect 3454 2418 3458 2422
rect 3438 2368 3442 2372
rect 3358 2358 3362 2362
rect 3382 2358 3386 2362
rect 3398 2358 3402 2362
rect 3462 2358 3466 2362
rect 3318 2338 3322 2342
rect 3246 2308 3250 2312
rect 3254 2308 3258 2312
rect 3198 2288 3202 2292
rect 3214 2288 3218 2292
rect 3190 2268 3194 2272
rect 3174 2248 3178 2252
rect 3190 2258 3194 2262
rect 3182 2238 3186 2242
rect 3174 2218 3178 2222
rect 3182 2218 3186 2222
rect 3166 2188 3170 2192
rect 3190 2178 3194 2182
rect 3086 2158 3090 2162
rect 3150 2158 3154 2162
rect 3214 2278 3218 2282
rect 3390 2338 3394 2342
rect 3414 2338 3418 2342
rect 3430 2338 3434 2342
rect 3326 2328 3330 2332
rect 3334 2328 3338 2332
rect 3350 2328 3354 2332
rect 3270 2318 3274 2322
rect 3310 2318 3314 2322
rect 3214 2248 3218 2252
rect 3222 2248 3226 2252
rect 3206 2238 3210 2242
rect 3238 2238 3242 2242
rect 3246 2218 3250 2222
rect 3262 2218 3266 2222
rect 3222 2208 3226 2212
rect 3334 2308 3338 2312
rect 3318 2288 3322 2292
rect 3350 2288 3354 2292
rect 3366 2328 3370 2332
rect 3382 2328 3386 2332
rect 3414 2318 3418 2322
rect 3446 2328 3450 2332
rect 3478 2338 3482 2342
rect 3390 2308 3394 2312
rect 3422 2308 3426 2312
rect 3454 2308 3458 2312
rect 3414 2298 3418 2302
rect 3374 2288 3378 2292
rect 3310 2268 3314 2272
rect 3286 2238 3290 2242
rect 3318 2238 3322 2242
rect 3398 2268 3402 2272
rect 3398 2248 3402 2252
rect 3342 2228 3346 2232
rect 3390 2218 3394 2222
rect 3326 2178 3330 2182
rect 3238 2168 3242 2172
rect 3310 2168 3314 2172
rect 3230 2158 3234 2162
rect 3294 2158 3298 2162
rect 3150 2148 3154 2152
rect 3190 2148 3194 2152
rect 3214 2148 3218 2152
rect 3230 2148 3234 2152
rect 3286 2148 3290 2152
rect 3070 2138 3074 2142
rect 3030 2118 3034 2122
rect 3042 2103 3046 2107
rect 3049 2103 3053 2107
rect 3054 2088 3058 2092
rect 3046 2078 3050 2082
rect 3038 2068 3042 2072
rect 3134 2128 3138 2132
rect 3166 2128 3170 2132
rect 3078 2118 3082 2122
rect 3078 2088 3082 2092
rect 3110 2088 3114 2092
rect 3070 2078 3074 2082
rect 3086 2078 3090 2082
rect 3102 2078 3106 2082
rect 3062 2068 3066 2072
rect 3070 2068 3074 2072
rect 3094 2068 3098 2072
rect 2982 2048 2986 2052
rect 3054 2048 3058 2052
rect 2998 2038 3002 2042
rect 3006 2038 3010 2042
rect 2966 2028 2970 2032
rect 2942 2018 2946 2022
rect 2958 2018 2962 2022
rect 2838 1988 2842 1992
rect 2862 1988 2866 1992
rect 2910 1988 2914 1992
rect 2774 1948 2778 1952
rect 2798 1948 2802 1952
rect 2822 1948 2826 1952
rect 2846 1948 2850 1952
rect 2766 1938 2770 1942
rect 2742 1918 2746 1922
rect 2750 1918 2754 1922
rect 2718 1888 2722 1892
rect 2710 1878 2714 1882
rect 2702 1868 2706 1872
rect 2734 1858 2738 1862
rect 2622 1848 2626 1852
rect 2598 1828 2602 1832
rect 2582 1818 2586 1822
rect 2598 1798 2602 1802
rect 2566 1778 2570 1782
rect 2534 1748 2538 1752
rect 2598 1748 2602 1752
rect 2590 1738 2594 1742
rect 2574 1728 2578 1732
rect 2510 1718 2514 1722
rect 2502 1708 2506 1712
rect 2486 1698 2490 1702
rect 2470 1668 2474 1672
rect 2398 1648 2402 1652
rect 2558 1708 2562 1712
rect 2542 1698 2546 1702
rect 2550 1688 2554 1692
rect 2542 1678 2546 1682
rect 2478 1658 2482 1662
rect 2494 1658 2498 1662
rect 2518 1658 2522 1662
rect 2550 1658 2554 1662
rect 2462 1648 2466 1652
rect 2574 1698 2578 1702
rect 2598 1698 2602 1702
rect 2582 1688 2586 1692
rect 2590 1678 2594 1682
rect 2582 1668 2586 1672
rect 2630 1808 2634 1812
rect 2638 1808 2642 1812
rect 2622 1718 2626 1722
rect 2622 1678 2626 1682
rect 2654 1798 2658 1802
rect 2670 1818 2674 1822
rect 2742 1848 2746 1852
rect 2758 1848 2762 1852
rect 2702 1828 2706 1832
rect 2710 1828 2714 1832
rect 2750 1828 2754 1832
rect 2678 1798 2682 1802
rect 2670 1778 2674 1782
rect 2662 1748 2666 1752
rect 2646 1728 2650 1732
rect 2694 1738 2698 1742
rect 2678 1708 2682 1712
rect 2686 1708 2690 1712
rect 2678 1678 2682 1682
rect 2686 1678 2690 1682
rect 2630 1668 2634 1672
rect 2582 1658 2586 1662
rect 2606 1658 2610 1662
rect 2654 1648 2658 1652
rect 2438 1628 2442 1632
rect 2454 1628 2458 1632
rect 2422 1608 2426 1612
rect 2422 1588 2426 1592
rect 2430 1588 2434 1592
rect 2454 1588 2458 1592
rect 2422 1568 2426 1572
rect 2414 1558 2418 1562
rect 2366 1498 2370 1502
rect 2454 1548 2458 1552
rect 2414 1538 2418 1542
rect 2446 1538 2450 1542
rect 2406 1528 2410 1532
rect 2574 1638 2578 1642
rect 2606 1638 2610 1642
rect 2638 1638 2642 1642
rect 2558 1628 2562 1632
rect 2486 1608 2490 1612
rect 2538 1603 2542 1607
rect 2545 1603 2549 1607
rect 2494 1588 2498 1592
rect 2510 1568 2514 1572
rect 2542 1568 2546 1572
rect 2630 1578 2634 1582
rect 2606 1568 2610 1572
rect 2550 1558 2554 1562
rect 2558 1558 2562 1562
rect 2358 1478 2362 1482
rect 2406 1478 2410 1482
rect 2366 1398 2370 1402
rect 2350 1388 2354 1392
rect 2342 1378 2346 1382
rect 2254 1348 2258 1352
rect 2262 1348 2266 1352
rect 2262 1298 2266 1302
rect 2214 1288 2218 1292
rect 2262 1278 2266 1282
rect 2206 1268 2210 1272
rect 2238 1268 2242 1272
rect 2190 1228 2194 1232
rect 2294 1328 2298 1332
rect 2302 1328 2306 1332
rect 2294 1288 2298 1292
rect 2286 1278 2290 1282
rect 2382 1398 2386 1402
rect 2374 1368 2378 1372
rect 2326 1348 2330 1352
rect 2358 1358 2362 1362
rect 2342 1348 2346 1352
rect 2318 1308 2322 1312
rect 2318 1278 2322 1282
rect 2446 1518 2450 1522
rect 2454 1518 2458 1522
rect 2486 1508 2490 1512
rect 2462 1478 2466 1482
rect 2478 1478 2482 1482
rect 2430 1468 2434 1472
rect 2406 1458 2410 1462
rect 2422 1458 2426 1462
rect 2414 1448 2418 1452
rect 2430 1448 2434 1452
rect 2414 1408 2418 1412
rect 2390 1348 2394 1352
rect 2406 1348 2410 1352
rect 2422 1348 2426 1352
rect 2382 1328 2386 1332
rect 2366 1308 2370 1312
rect 2374 1308 2378 1312
rect 2454 1448 2458 1452
rect 2470 1438 2474 1442
rect 2478 1358 2482 1362
rect 2390 1298 2394 1302
rect 2430 1298 2434 1302
rect 2382 1288 2386 1292
rect 2406 1288 2410 1292
rect 2438 1288 2442 1292
rect 2462 1288 2466 1292
rect 2526 1528 2530 1532
rect 2518 1518 2522 1522
rect 2534 1498 2538 1502
rect 2558 1548 2562 1552
rect 2574 1548 2578 1552
rect 2654 1558 2658 1562
rect 2678 1638 2682 1642
rect 2694 1608 2698 1612
rect 2694 1598 2698 1602
rect 2678 1588 2682 1592
rect 2662 1548 2666 1552
rect 2582 1538 2586 1542
rect 2598 1538 2602 1542
rect 2686 1538 2690 1542
rect 2598 1528 2602 1532
rect 2622 1528 2626 1532
rect 2638 1528 2642 1532
rect 2558 1498 2562 1502
rect 2582 1498 2586 1502
rect 2590 1498 2594 1502
rect 2582 1478 2586 1482
rect 2510 1458 2514 1462
rect 2558 1438 2562 1442
rect 2510 1408 2514 1412
rect 2558 1408 2562 1412
rect 2538 1403 2542 1407
rect 2545 1403 2549 1407
rect 2510 1398 2514 1402
rect 2502 1388 2506 1392
rect 2526 1368 2530 1372
rect 2494 1358 2498 1362
rect 2510 1348 2514 1352
rect 2542 1358 2546 1362
rect 2502 1328 2506 1332
rect 2486 1318 2490 1322
rect 2478 1308 2482 1312
rect 2382 1278 2386 1282
rect 2470 1278 2474 1282
rect 2518 1288 2522 1292
rect 2606 1468 2610 1472
rect 2598 1458 2602 1462
rect 2638 1498 2642 1502
rect 2630 1488 2634 1492
rect 2638 1398 2642 1402
rect 2614 1388 2618 1392
rect 2598 1358 2602 1362
rect 2614 1358 2618 1362
rect 2622 1358 2626 1362
rect 2574 1348 2578 1352
rect 2670 1528 2674 1532
rect 2662 1518 2666 1522
rect 2678 1498 2682 1502
rect 2686 1488 2690 1492
rect 2670 1478 2674 1482
rect 2662 1468 2666 1472
rect 2678 1458 2682 1462
rect 2670 1448 2674 1452
rect 2686 1448 2690 1452
rect 2670 1388 2674 1392
rect 2598 1338 2602 1342
rect 2638 1338 2642 1342
rect 2566 1328 2570 1332
rect 2574 1328 2578 1332
rect 2582 1328 2586 1332
rect 2582 1308 2586 1312
rect 2526 1278 2530 1282
rect 2534 1278 2538 1282
rect 2270 1258 2274 1262
rect 2286 1258 2290 1262
rect 2230 1248 2234 1252
rect 2230 1218 2234 1222
rect 2206 1198 2210 1202
rect 2214 1198 2218 1202
rect 2174 1158 2178 1162
rect 2294 1228 2298 1232
rect 2270 1218 2274 1222
rect 2238 1188 2242 1192
rect 2198 1148 2202 1152
rect 2214 1148 2218 1152
rect 2230 1148 2234 1152
rect 2262 1148 2266 1152
rect 2270 1148 2274 1152
rect 2174 1138 2178 1142
rect 2158 1058 2162 1062
rect 2142 998 2146 1002
rect 2254 1138 2258 1142
rect 2206 1128 2210 1132
rect 2182 1088 2186 1092
rect 2238 1128 2242 1132
rect 2182 1078 2186 1082
rect 2230 1078 2234 1082
rect 2246 1098 2250 1102
rect 2214 1068 2218 1072
rect 2174 1048 2178 1052
rect 2166 1038 2170 1042
rect 2230 1038 2234 1042
rect 2182 968 2186 972
rect 2190 958 2194 962
rect 2254 988 2258 992
rect 2222 968 2226 972
rect 2230 968 2234 972
rect 2158 948 2162 952
rect 2198 948 2202 952
rect 2222 948 2226 952
rect 2302 1218 2306 1222
rect 2326 1248 2330 1252
rect 2326 1228 2330 1232
rect 2326 1218 2330 1222
rect 2294 1088 2298 1092
rect 2318 1158 2322 1162
rect 2318 1118 2322 1122
rect 2310 1098 2314 1102
rect 2302 1078 2306 1082
rect 2350 1248 2354 1252
rect 2374 1178 2378 1182
rect 2334 1168 2338 1172
rect 2366 1148 2370 1152
rect 2366 1118 2370 1122
rect 2350 1098 2354 1102
rect 2350 1088 2354 1092
rect 2366 1078 2370 1082
rect 2382 1078 2386 1082
rect 2286 1058 2290 1062
rect 2318 1058 2322 1062
rect 2334 1058 2338 1062
rect 2278 1048 2282 1052
rect 2286 1048 2290 1052
rect 2310 1048 2314 1052
rect 2326 1048 2330 1052
rect 2302 1038 2306 1042
rect 2310 1038 2314 1042
rect 2278 1008 2282 1012
rect 2270 998 2274 1002
rect 2150 938 2154 942
rect 2182 938 2186 942
rect 2222 938 2226 942
rect 2262 938 2266 942
rect 2134 928 2138 932
rect 2150 898 2154 902
rect 2174 898 2178 902
rect 2134 888 2138 892
rect 2126 868 2130 872
rect 2158 868 2162 872
rect 2198 898 2202 902
rect 2198 888 2202 892
rect 2102 858 2106 862
rect 2110 838 2114 842
rect 2094 808 2098 812
rect 2110 808 2114 812
rect 2062 768 2066 772
rect 1990 758 1994 762
rect 2046 758 2050 762
rect 2070 758 2074 762
rect 1950 738 1954 742
rect 1990 738 1994 742
rect 1934 728 1938 732
rect 1958 728 1962 732
rect 1974 728 1978 732
rect 2030 748 2034 752
rect 2086 748 2090 752
rect 2014 728 2018 732
rect 2062 728 2066 732
rect 2102 728 2106 732
rect 1998 718 2002 722
rect 2054 718 2058 722
rect 1942 708 1946 712
rect 1950 678 1954 682
rect 2006 678 2010 682
rect 2102 708 2106 712
rect 2026 703 2030 707
rect 2033 703 2037 707
rect 2126 848 2130 852
rect 2206 868 2210 872
rect 2230 878 2234 882
rect 2142 858 2146 862
rect 2150 858 2154 862
rect 2134 838 2138 842
rect 2150 798 2154 802
rect 2206 788 2210 792
rect 2150 758 2154 762
rect 2166 758 2170 762
rect 2118 748 2122 752
rect 2126 748 2130 752
rect 2126 728 2130 732
rect 2134 718 2138 722
rect 2078 678 2082 682
rect 2014 668 2018 672
rect 2022 668 2026 672
rect 1910 658 1914 662
rect 2014 658 2018 662
rect 2054 658 2058 662
rect 2078 658 2082 662
rect 1886 638 1890 642
rect 1918 638 1922 642
rect 1942 638 1946 642
rect 1798 568 1802 572
rect 1862 568 1866 572
rect 1774 558 1778 562
rect 1814 558 1818 562
rect 1838 558 1842 562
rect 1686 548 1690 552
rect 1766 548 1770 552
rect 1710 538 1714 542
rect 1686 528 1690 532
rect 1670 518 1674 522
rect 1710 518 1714 522
rect 1678 488 1682 492
rect 1582 468 1586 472
rect 1598 468 1602 472
rect 1614 468 1618 472
rect 1646 468 1650 472
rect 1614 458 1618 462
rect 1638 458 1642 462
rect 1582 438 1586 442
rect 1622 418 1626 422
rect 1638 418 1642 422
rect 1630 378 1634 382
rect 1566 368 1570 372
rect 1614 348 1618 352
rect 1622 348 1626 352
rect 1582 308 1586 312
rect 1542 298 1546 302
rect 1614 328 1618 332
rect 1550 278 1554 282
rect 1582 278 1586 282
rect 1598 278 1602 282
rect 1614 278 1618 282
rect 1542 268 1546 272
rect 1566 268 1570 272
rect 1566 248 1570 252
rect 1534 238 1538 242
rect 1598 258 1602 262
rect 1606 258 1610 262
rect 1606 238 1610 242
rect 1526 218 1530 222
rect 1582 218 1586 222
rect 1486 148 1490 152
rect 1514 203 1518 207
rect 1521 203 1525 207
rect 1662 448 1666 452
rect 1686 448 1690 452
rect 1670 438 1674 442
rect 1654 418 1658 422
rect 1694 418 1698 422
rect 1678 378 1682 382
rect 1670 368 1674 372
rect 1646 358 1650 362
rect 1678 348 1682 352
rect 1694 348 1698 352
rect 1670 318 1674 322
rect 1662 308 1666 312
rect 1646 278 1650 282
rect 1798 518 1802 522
rect 1790 508 1794 512
rect 1750 488 1754 492
rect 1758 458 1762 462
rect 1774 458 1778 462
rect 1822 498 1826 502
rect 1830 488 1834 492
rect 1870 548 1874 552
rect 1862 518 1866 522
rect 1878 518 1882 522
rect 1934 598 1938 602
rect 1918 558 1922 562
rect 1902 548 1906 552
rect 1926 548 1930 552
rect 2046 648 2050 652
rect 2126 658 2130 662
rect 2158 748 2162 752
rect 2190 748 2194 752
rect 2230 848 2234 852
rect 2286 978 2290 982
rect 2270 868 2274 872
rect 2294 918 2298 922
rect 2302 908 2306 912
rect 2334 968 2338 972
rect 2358 968 2362 972
rect 2374 1058 2378 1062
rect 2422 1258 2426 1262
rect 2438 1258 2442 1262
rect 2462 1258 2466 1262
rect 2478 1258 2482 1262
rect 2494 1268 2498 1272
rect 2494 1258 2498 1262
rect 2486 1238 2490 1242
rect 2430 1218 2434 1222
rect 2494 1218 2498 1222
rect 2414 1188 2418 1192
rect 2446 1208 2450 1212
rect 2590 1258 2594 1262
rect 2550 1248 2554 1252
rect 2574 1248 2578 1252
rect 2558 1238 2562 1242
rect 2538 1203 2542 1207
rect 2545 1203 2549 1207
rect 2526 1198 2530 1202
rect 2566 1218 2570 1222
rect 2430 1178 2434 1182
rect 2446 1178 2450 1182
rect 2406 1158 2410 1162
rect 2414 1158 2418 1162
rect 2502 1168 2506 1172
rect 2398 1138 2402 1142
rect 2510 1138 2514 1142
rect 2518 1138 2522 1142
rect 2454 1128 2458 1132
rect 2486 1128 2490 1132
rect 2526 1128 2530 1132
rect 2550 1128 2554 1132
rect 2430 1088 2434 1092
rect 2486 1108 2490 1112
rect 2414 1058 2418 1062
rect 2430 1058 2434 1062
rect 2398 1048 2402 1052
rect 2446 1028 2450 1032
rect 2406 1008 2410 1012
rect 2390 988 2394 992
rect 2366 958 2370 962
rect 2382 958 2386 962
rect 2326 948 2330 952
rect 2374 948 2378 952
rect 2334 938 2338 942
rect 2302 878 2306 882
rect 2342 898 2346 902
rect 2310 868 2314 872
rect 2414 938 2418 942
rect 2366 908 2370 912
rect 2350 878 2354 882
rect 2342 858 2346 862
rect 2294 848 2298 852
rect 2326 848 2330 852
rect 2262 838 2266 842
rect 2254 808 2258 812
rect 2222 758 2226 762
rect 2294 758 2298 762
rect 2342 758 2346 762
rect 2278 748 2282 752
rect 2310 748 2314 752
rect 2214 738 2218 742
rect 2222 738 2226 742
rect 2246 738 2250 742
rect 2286 738 2290 742
rect 2174 718 2178 722
rect 2166 688 2170 692
rect 2278 718 2282 722
rect 2262 708 2266 712
rect 2310 708 2314 712
rect 2334 708 2338 712
rect 2222 688 2226 692
rect 2182 678 2186 682
rect 2214 678 2218 682
rect 2150 668 2154 672
rect 2094 648 2098 652
rect 2190 668 2194 672
rect 2198 658 2202 662
rect 2070 638 2074 642
rect 2086 638 2090 642
rect 2134 638 2138 642
rect 2166 638 2170 642
rect 2174 618 2178 622
rect 1982 598 1986 602
rect 2110 598 2114 602
rect 1998 578 2002 582
rect 2110 578 2114 582
rect 1998 558 2002 562
rect 1910 538 1914 542
rect 1950 538 1954 542
rect 1966 538 1970 542
rect 2070 558 2074 562
rect 2118 558 2122 562
rect 1998 548 2002 552
rect 2046 548 2050 552
rect 1998 538 2002 542
rect 2006 538 2010 542
rect 1894 498 1898 502
rect 1870 478 1874 482
rect 1886 478 1890 482
rect 1894 478 1898 482
rect 1830 468 1834 472
rect 1790 448 1794 452
rect 1726 398 1730 402
rect 1742 438 1746 442
rect 1782 438 1786 442
rect 1718 388 1722 392
rect 1814 448 1818 452
rect 1822 438 1826 442
rect 1806 428 1810 432
rect 1750 368 1754 372
rect 1734 348 1738 352
rect 1758 348 1762 352
rect 1710 328 1714 332
rect 1686 318 1690 322
rect 1726 308 1730 312
rect 1702 288 1706 292
rect 1686 278 1690 282
rect 1710 278 1714 282
rect 1774 398 1778 402
rect 1790 358 1794 362
rect 1774 348 1778 352
rect 1806 348 1810 352
rect 1822 348 1826 352
rect 1806 328 1810 332
rect 1790 318 1794 322
rect 1766 278 1770 282
rect 1814 308 1818 312
rect 1862 458 1866 462
rect 1846 438 1850 442
rect 1854 388 1858 392
rect 1846 358 1850 362
rect 1838 348 1842 352
rect 1878 448 1882 452
rect 1870 428 1874 432
rect 1838 308 1842 312
rect 1630 258 1634 262
rect 1646 258 1650 262
rect 1718 258 1722 262
rect 1742 258 1746 262
rect 1766 258 1770 262
rect 1790 258 1794 262
rect 1630 248 1634 252
rect 1646 248 1650 252
rect 1678 248 1682 252
rect 1622 228 1626 232
rect 1654 238 1658 242
rect 1542 158 1546 162
rect 1558 158 1562 162
rect 1590 158 1594 162
rect 1638 158 1642 162
rect 1534 148 1538 152
rect 1542 148 1546 152
rect 1494 138 1498 142
rect 1526 128 1530 132
rect 1486 118 1490 122
rect 1534 98 1538 102
rect 1398 78 1402 82
rect 1414 78 1418 82
rect 1446 78 1450 82
rect 1462 78 1466 82
rect 1502 78 1506 82
rect 1286 68 1290 72
rect 1278 58 1282 62
rect 1318 58 1322 62
rect 1102 28 1106 32
rect 1214 8 1218 12
rect 1270 8 1274 12
rect 1350 58 1354 62
rect 1374 58 1378 62
rect 1430 68 1434 72
rect 1422 58 1426 62
rect 1438 58 1442 62
rect 1470 68 1474 72
rect 1486 68 1490 72
rect 1518 68 1522 72
rect 1558 138 1562 142
rect 1590 138 1594 142
rect 1598 138 1602 142
rect 1558 128 1562 132
rect 1590 128 1594 132
rect 1550 118 1554 122
rect 1614 118 1618 122
rect 1638 98 1642 102
rect 1558 78 1562 82
rect 1614 78 1618 82
rect 1478 58 1482 62
rect 1526 58 1530 62
rect 1406 48 1410 52
rect 1438 48 1442 52
rect 1566 38 1570 42
rect 1566 18 1570 22
rect 1622 48 1626 52
rect 1638 48 1642 52
rect 1662 228 1666 232
rect 1678 218 1682 222
rect 1678 158 1682 162
rect 1670 148 1674 152
rect 1654 138 1658 142
rect 1662 138 1666 142
rect 1726 198 1730 202
rect 1694 148 1698 152
rect 1702 148 1706 152
rect 1702 128 1706 132
rect 1726 118 1730 122
rect 1670 98 1674 102
rect 1774 248 1778 252
rect 1806 248 1810 252
rect 1822 248 1826 252
rect 1878 378 1882 382
rect 1926 518 1930 522
rect 1910 458 1914 462
rect 1902 448 1906 452
rect 1910 448 1914 452
rect 1934 498 1938 502
rect 1990 518 1994 522
rect 1974 508 1978 512
rect 1982 498 1986 502
rect 2062 528 2066 532
rect 2094 528 2098 532
rect 2054 518 2058 522
rect 2026 503 2030 507
rect 2033 503 2037 507
rect 2014 488 2018 492
rect 2030 478 2034 482
rect 2046 478 2050 482
rect 2062 478 2066 482
rect 2086 478 2090 482
rect 1950 458 1954 462
rect 1990 468 1994 472
rect 2006 468 2010 472
rect 2022 468 2026 472
rect 1966 458 1970 462
rect 1918 428 1922 432
rect 1926 408 1930 412
rect 1918 398 1922 402
rect 1894 378 1898 382
rect 1902 368 1906 372
rect 1894 348 1898 352
rect 1942 378 1946 382
rect 1974 438 1978 442
rect 1950 368 1954 372
rect 1990 458 1994 462
rect 2022 418 2026 422
rect 2006 378 2010 382
rect 1950 358 1954 362
rect 1982 358 1986 362
rect 1990 358 1994 362
rect 2054 458 2058 462
rect 2070 458 2074 462
rect 2078 448 2082 452
rect 2094 428 2098 432
rect 2054 418 2058 422
rect 1950 348 1954 352
rect 1974 348 1978 352
rect 2022 348 2026 352
rect 1998 338 2002 342
rect 2006 338 2010 342
rect 1886 328 1890 332
rect 1910 328 1914 332
rect 1862 308 1866 312
rect 1854 298 1858 302
rect 1854 288 1858 292
rect 1862 288 1866 292
rect 1862 268 1866 272
rect 1886 268 1890 272
rect 1870 248 1874 252
rect 1910 308 1914 312
rect 1902 298 1906 302
rect 1942 298 1946 302
rect 2022 328 2026 332
rect 2046 318 2050 322
rect 1998 298 2002 302
rect 1910 268 1914 272
rect 1886 248 1890 252
rect 1902 248 1906 252
rect 2026 303 2030 307
rect 2033 303 2037 307
rect 1926 248 1930 252
rect 1846 238 1850 242
rect 1878 238 1882 242
rect 1910 238 1914 242
rect 1958 238 1962 242
rect 1846 228 1850 232
rect 1878 228 1882 232
rect 1838 198 1842 202
rect 1862 208 1866 212
rect 1870 198 1874 202
rect 1742 158 1746 162
rect 1758 148 1762 152
rect 1814 148 1818 152
rect 1766 128 1770 132
rect 1766 108 1770 112
rect 1782 108 1786 112
rect 1814 108 1818 112
rect 1734 98 1738 102
rect 1766 98 1770 102
rect 1686 78 1690 82
rect 1694 78 1698 82
rect 1686 58 1690 62
rect 1742 58 1746 62
rect 1814 98 1818 102
rect 1862 138 1866 142
rect 1854 128 1858 132
rect 1830 108 1834 112
rect 1822 58 1826 62
rect 1782 48 1786 52
rect 1702 38 1706 42
rect 1774 38 1778 42
rect 1646 18 1650 22
rect 1486 8 1490 12
rect 1542 8 1546 12
rect 1598 8 1602 12
rect 1614 8 1618 12
rect 1514 3 1518 7
rect 1521 3 1525 7
rect 1814 48 1818 52
rect 1974 228 1978 232
rect 1982 228 1986 232
rect 1990 228 1994 232
rect 1942 208 1946 212
rect 1910 178 1914 182
rect 1910 158 1914 162
rect 1942 158 1946 162
rect 1950 148 1954 152
rect 2006 148 2010 152
rect 2070 358 2074 362
rect 2070 348 2074 352
rect 2214 658 2218 662
rect 2166 578 2170 582
rect 2206 578 2210 582
rect 2150 558 2154 562
rect 2158 558 2162 562
rect 2150 548 2154 552
rect 2254 648 2258 652
rect 2198 538 2202 542
rect 2382 898 2386 902
rect 2390 888 2394 892
rect 2414 858 2418 862
rect 2374 848 2378 852
rect 2406 798 2410 802
rect 2430 988 2434 992
rect 2478 1018 2482 1022
rect 2446 948 2450 952
rect 2526 1098 2530 1102
rect 2558 1098 2562 1102
rect 2494 1088 2498 1092
rect 2542 1068 2546 1072
rect 2622 1328 2626 1332
rect 2654 1328 2658 1332
rect 2646 1318 2650 1322
rect 2606 1308 2610 1312
rect 2606 1298 2610 1302
rect 2854 1938 2858 1942
rect 2870 1938 2874 1942
rect 2814 1928 2818 1932
rect 2774 1918 2778 1922
rect 2790 1918 2794 1922
rect 2774 1868 2778 1872
rect 2854 1908 2858 1912
rect 2838 1888 2842 1892
rect 3054 2008 3058 2012
rect 2990 1998 2994 2002
rect 2974 1988 2978 1992
rect 2966 1978 2970 1982
rect 2950 1968 2954 1972
rect 2918 1958 2922 1962
rect 2958 1958 2962 1962
rect 2926 1948 2930 1952
rect 2918 1938 2922 1942
rect 2942 1938 2946 1942
rect 2878 1928 2882 1932
rect 2910 1908 2914 1912
rect 3014 1968 3018 1972
rect 3030 1968 3034 1972
rect 3006 1948 3010 1952
rect 2982 1928 2986 1932
rect 2966 1908 2970 1912
rect 3046 1938 3050 1942
rect 3014 1908 3018 1912
rect 2990 1898 2994 1902
rect 3042 1903 3046 1907
rect 3049 1903 3053 1907
rect 3134 2068 3138 2072
rect 3182 2088 3186 2092
rect 3150 2078 3154 2082
rect 3198 2078 3202 2082
rect 3214 2098 3218 2102
rect 3078 2048 3082 2052
rect 3182 2048 3186 2052
rect 3070 1968 3074 1972
rect 3070 1938 3074 1942
rect 3126 2028 3130 2032
rect 3142 2018 3146 2022
rect 3086 2008 3090 2012
rect 3110 1998 3114 2002
rect 3022 1898 3026 1902
rect 3062 1898 3066 1902
rect 2870 1888 2874 1892
rect 2894 1888 2898 1892
rect 2926 1888 2930 1892
rect 3102 1938 3106 1942
rect 3118 1988 3122 1992
rect 3134 1988 3138 1992
rect 3126 1968 3130 1972
rect 3222 2048 3226 2052
rect 3206 2038 3210 2042
rect 3198 1998 3202 2002
rect 3150 1978 3154 1982
rect 3174 1978 3178 1982
rect 3142 1958 3146 1962
rect 3158 1958 3162 1962
rect 3190 1958 3194 1962
rect 3334 2148 3338 2152
rect 3374 2148 3378 2152
rect 3270 2138 3274 2142
rect 3262 2118 3266 2122
rect 3262 2088 3266 2092
rect 3286 2128 3290 2132
rect 3350 2128 3354 2132
rect 3302 2108 3306 2112
rect 3326 2108 3330 2112
rect 3382 2118 3386 2122
rect 3358 2098 3362 2102
rect 3510 2458 3514 2462
rect 3518 2458 3522 2462
rect 3534 2448 3538 2452
rect 3494 2348 3498 2352
rect 3502 2348 3506 2352
rect 3454 2268 3458 2272
rect 3446 2248 3450 2252
rect 3510 2248 3514 2252
rect 3422 2218 3426 2222
rect 3422 2208 3426 2212
rect 3470 2238 3474 2242
rect 3430 2198 3434 2202
rect 3478 2198 3482 2202
rect 3438 2188 3442 2192
rect 3430 2158 3434 2162
rect 3406 2128 3410 2132
rect 3454 2128 3458 2132
rect 3390 2098 3394 2102
rect 3366 2078 3370 2082
rect 3326 2068 3330 2072
rect 3350 2068 3354 2072
rect 3374 2068 3378 2072
rect 3318 2058 3322 2062
rect 3366 2058 3370 2062
rect 3350 2048 3354 2052
rect 3294 2038 3298 2042
rect 3238 2008 3242 2012
rect 3230 1988 3234 1992
rect 3190 1948 3194 1952
rect 3206 1948 3210 1952
rect 3246 1968 3250 1972
rect 3294 1968 3298 1972
rect 3270 1958 3274 1962
rect 3262 1948 3266 1952
rect 3278 1948 3282 1952
rect 3302 1958 3306 1962
rect 3358 1958 3362 1962
rect 3206 1938 3210 1942
rect 3230 1938 3234 1942
rect 3302 1938 3306 1942
rect 3158 1928 3162 1932
rect 3238 1928 3242 1932
rect 3118 1908 3122 1912
rect 3142 1888 3146 1892
rect 2846 1878 2850 1882
rect 3118 1878 3122 1882
rect 2830 1868 2834 1872
rect 2870 1868 2874 1872
rect 2846 1858 2850 1862
rect 2822 1848 2826 1852
rect 2790 1828 2794 1832
rect 2814 1828 2818 1832
rect 2854 1828 2858 1832
rect 2766 1808 2770 1812
rect 2758 1798 2762 1802
rect 2790 1798 2794 1802
rect 2798 1788 2802 1792
rect 2718 1778 2722 1782
rect 2726 1768 2730 1772
rect 2790 1768 2794 1772
rect 2830 1758 2834 1762
rect 2718 1748 2722 1752
rect 2750 1748 2754 1752
rect 2806 1748 2810 1752
rect 2726 1738 2730 1742
rect 2838 1738 2842 1742
rect 2902 1868 2906 1872
rect 2926 1868 2930 1872
rect 2998 1868 3002 1872
rect 3086 1868 3090 1872
rect 2942 1858 2946 1862
rect 2990 1858 2994 1862
rect 3006 1858 3010 1862
rect 3078 1858 3082 1862
rect 2958 1848 2962 1852
rect 2902 1818 2906 1822
rect 2878 1798 2882 1802
rect 2934 1808 2938 1812
rect 2918 1768 2922 1772
rect 2998 1848 3002 1852
rect 3038 1848 3042 1852
rect 2998 1838 3002 1842
rect 2942 1778 2946 1782
rect 2894 1748 2898 1752
rect 2886 1738 2890 1742
rect 2814 1728 2818 1732
rect 2710 1708 2714 1712
rect 2774 1708 2778 1712
rect 2742 1698 2746 1702
rect 2782 1698 2786 1702
rect 2710 1688 2714 1692
rect 2718 1678 2722 1682
rect 2726 1668 2730 1672
rect 2782 1668 2786 1672
rect 2750 1658 2754 1662
rect 2766 1658 2770 1662
rect 2734 1648 2738 1652
rect 2774 1628 2778 1632
rect 2710 1548 2714 1552
rect 2718 1508 2722 1512
rect 2750 1608 2754 1612
rect 2822 1678 2826 1682
rect 2814 1658 2818 1662
rect 2846 1658 2850 1662
rect 2830 1638 2834 1642
rect 2798 1598 2802 1602
rect 2798 1588 2802 1592
rect 2734 1568 2738 1572
rect 2734 1558 2738 1562
rect 2750 1558 2754 1562
rect 2806 1578 2810 1582
rect 2894 1638 2898 1642
rect 2878 1628 2882 1632
rect 2854 1578 2858 1582
rect 2838 1568 2842 1572
rect 2830 1558 2834 1562
rect 2910 1718 2914 1722
rect 2910 1668 2914 1672
rect 2966 1748 2970 1752
rect 3230 1898 3234 1902
rect 3222 1878 3226 1882
rect 3318 1928 3322 1932
rect 3326 1888 3330 1892
rect 3318 1878 3322 1882
rect 3150 1868 3154 1872
rect 3102 1858 3106 1862
rect 3118 1858 3122 1862
rect 3102 1818 3106 1822
rect 3094 1808 3098 1812
rect 3030 1758 3034 1762
rect 3086 1758 3090 1762
rect 3062 1748 3066 1752
rect 2942 1738 2946 1742
rect 3070 1738 3074 1742
rect 3086 1738 3090 1742
rect 2950 1718 2954 1722
rect 2998 1728 3002 1732
rect 2974 1718 2978 1722
rect 2966 1688 2970 1692
rect 2934 1668 2938 1672
rect 2926 1648 2930 1652
rect 2918 1628 2922 1632
rect 2902 1588 2906 1592
rect 2870 1568 2874 1572
rect 2878 1568 2882 1572
rect 2894 1568 2898 1572
rect 2846 1548 2850 1552
rect 2862 1548 2866 1552
rect 2878 1548 2882 1552
rect 2790 1528 2794 1532
rect 2734 1518 2738 1522
rect 2806 1518 2810 1522
rect 2758 1508 2762 1512
rect 2726 1498 2730 1502
rect 2726 1488 2730 1492
rect 2710 1468 2714 1472
rect 2734 1468 2738 1472
rect 2798 1468 2802 1472
rect 2758 1458 2762 1462
rect 2774 1458 2778 1462
rect 2718 1448 2722 1452
rect 2774 1448 2778 1452
rect 2822 1528 2826 1532
rect 2862 1528 2866 1532
rect 2942 1648 2946 1652
rect 2958 1648 2962 1652
rect 2950 1558 2954 1562
rect 2982 1678 2986 1682
rect 3078 1708 3082 1712
rect 3042 1703 3046 1707
rect 3049 1703 3053 1707
rect 3094 1698 3098 1702
rect 3006 1688 3010 1692
rect 3062 1688 3066 1692
rect 3158 1848 3162 1852
rect 3206 1858 3210 1862
rect 3222 1858 3226 1862
rect 3230 1858 3234 1862
rect 3174 1838 3178 1842
rect 3262 1858 3266 1862
rect 3254 1848 3258 1852
rect 3462 2068 3466 2072
rect 3430 2048 3434 2052
rect 3398 2018 3402 2022
rect 3430 1968 3434 1972
rect 3390 1958 3394 1962
rect 3414 1958 3418 1962
rect 3470 2008 3474 2012
rect 3558 2348 3562 2352
rect 3526 2298 3530 2302
rect 3550 2298 3554 2302
rect 3558 2298 3562 2302
rect 3558 2268 3562 2272
rect 3542 2248 3546 2252
rect 3542 2058 3546 2062
rect 3494 2018 3498 2022
rect 3486 1988 3490 1992
rect 3470 1968 3474 1972
rect 3486 1968 3490 1972
rect 3446 1948 3450 1952
rect 3478 1948 3482 1952
rect 3382 1928 3386 1932
rect 3374 1888 3378 1892
rect 3454 1938 3458 1942
rect 3558 2048 3562 2052
rect 3526 2018 3530 2022
rect 3502 2008 3506 2012
rect 3502 1958 3506 1962
rect 3518 1978 3522 1982
rect 3518 1948 3522 1952
rect 3558 1948 3562 1952
rect 3518 1938 3522 1942
rect 3510 1898 3514 1902
rect 3478 1888 3482 1892
rect 3510 1878 3514 1882
rect 3526 1878 3530 1882
rect 3398 1868 3402 1872
rect 3454 1868 3458 1872
rect 3286 1848 3290 1852
rect 3150 1818 3154 1822
rect 3246 1818 3250 1822
rect 3278 1818 3282 1822
rect 3110 1758 3114 1762
rect 3230 1788 3234 1792
rect 3294 1788 3298 1792
rect 3286 1778 3290 1782
rect 3358 1778 3362 1782
rect 3366 1778 3370 1782
rect 3182 1758 3186 1762
rect 3262 1758 3266 1762
rect 3302 1758 3306 1762
rect 3406 1858 3410 1862
rect 3454 1859 3458 1863
rect 3398 1848 3402 1852
rect 3406 1848 3410 1852
rect 3558 1848 3562 1852
rect 3510 1828 3514 1832
rect 3438 1818 3442 1822
rect 3406 1778 3410 1782
rect 3110 1728 3114 1732
rect 3134 1728 3138 1732
rect 3206 1748 3210 1752
rect 3254 1748 3258 1752
rect 3358 1748 3362 1752
rect 3374 1748 3378 1752
rect 3230 1738 3234 1742
rect 3238 1738 3242 1742
rect 3262 1738 3266 1742
rect 3294 1738 3298 1742
rect 3350 1738 3354 1742
rect 3150 1728 3154 1732
rect 3206 1728 3210 1732
rect 3286 1728 3290 1732
rect 3142 1708 3146 1712
rect 3158 1688 3162 1692
rect 3174 1688 3178 1692
rect 3030 1678 3034 1682
rect 3030 1658 3034 1662
rect 3070 1658 3074 1662
rect 3102 1658 3106 1662
rect 3142 1658 3146 1662
rect 2990 1598 2994 1602
rect 2998 1588 3002 1592
rect 2974 1578 2978 1582
rect 2990 1568 2994 1572
rect 2934 1538 2938 1542
rect 2942 1538 2946 1542
rect 2910 1528 2914 1532
rect 2926 1518 2930 1522
rect 2942 1518 2946 1522
rect 2918 1508 2922 1512
rect 2934 1508 2938 1512
rect 2822 1488 2826 1492
rect 2886 1488 2890 1492
rect 2902 1488 2906 1492
rect 2846 1478 2850 1482
rect 2862 1478 2866 1482
rect 2886 1478 2890 1482
rect 2870 1468 2874 1472
rect 2830 1458 2834 1462
rect 2846 1458 2850 1462
rect 2814 1418 2818 1422
rect 2702 1388 2706 1392
rect 2862 1418 2866 1422
rect 2862 1398 2866 1402
rect 2838 1388 2842 1392
rect 2726 1368 2730 1372
rect 2782 1368 2786 1372
rect 2702 1358 2706 1362
rect 2766 1358 2770 1362
rect 2790 1358 2794 1362
rect 2838 1358 2842 1362
rect 2686 1348 2690 1352
rect 2726 1348 2730 1352
rect 2758 1348 2762 1352
rect 2678 1338 2682 1342
rect 2686 1328 2690 1332
rect 2710 1328 2714 1332
rect 2622 1268 2626 1272
rect 2646 1268 2650 1272
rect 2702 1268 2706 1272
rect 2614 1248 2618 1252
rect 2598 1228 2602 1232
rect 2606 1228 2610 1232
rect 2582 1178 2586 1182
rect 2574 1168 2578 1172
rect 2582 1168 2586 1172
rect 2638 1248 2642 1252
rect 2654 1248 2658 1252
rect 2630 1208 2634 1212
rect 2630 1198 2634 1202
rect 2614 1168 2618 1172
rect 2574 1138 2578 1142
rect 2538 1003 2542 1007
rect 2545 1003 2549 1007
rect 2558 968 2562 972
rect 2622 1078 2626 1082
rect 2638 1178 2642 1182
rect 2678 1158 2682 1162
rect 2734 1338 2738 1342
rect 2750 1338 2754 1342
rect 2718 1318 2722 1322
rect 2782 1308 2786 1312
rect 2910 1468 2914 1472
rect 2926 1468 2930 1472
rect 2886 1458 2890 1462
rect 2974 1518 2978 1522
rect 2950 1508 2954 1512
rect 2950 1498 2954 1502
rect 2942 1488 2946 1492
rect 2966 1478 2970 1482
rect 2974 1478 2978 1482
rect 3198 1708 3202 1712
rect 3214 1688 3218 1692
rect 3246 1678 3250 1682
rect 3262 1678 3266 1682
rect 3054 1648 3058 1652
rect 3086 1648 3090 1652
rect 3134 1648 3138 1652
rect 3174 1648 3178 1652
rect 3190 1648 3194 1652
rect 3254 1668 3258 1672
rect 3270 1668 3274 1672
rect 3206 1658 3210 1662
rect 3150 1638 3154 1642
rect 3198 1638 3202 1642
rect 3206 1638 3210 1642
rect 3118 1618 3122 1622
rect 3086 1608 3090 1612
rect 3134 1608 3138 1612
rect 3078 1558 3082 1562
rect 3006 1548 3010 1552
rect 3070 1548 3074 1552
rect 2990 1538 2994 1542
rect 3070 1538 3074 1542
rect 2998 1518 3002 1522
rect 3030 1518 3034 1522
rect 2990 1488 2994 1492
rect 3042 1503 3046 1507
rect 3049 1503 3053 1507
rect 3022 1498 3026 1502
rect 3006 1478 3010 1482
rect 3022 1478 3026 1482
rect 3030 1468 3034 1472
rect 3054 1468 3058 1472
rect 2974 1458 2978 1462
rect 2958 1448 2962 1452
rect 3030 1448 3034 1452
rect 3062 1448 3066 1452
rect 3062 1438 3066 1442
rect 2934 1428 2938 1432
rect 2990 1428 2994 1432
rect 2910 1408 2914 1412
rect 2886 1378 2890 1382
rect 2926 1358 2930 1362
rect 2814 1348 2818 1352
rect 2822 1348 2826 1352
rect 2862 1348 2866 1352
rect 2998 1378 3002 1382
rect 2942 1358 2946 1362
rect 2982 1358 2986 1362
rect 2958 1348 2962 1352
rect 2982 1348 2986 1352
rect 2998 1348 3002 1352
rect 2798 1338 2802 1342
rect 2814 1338 2818 1342
rect 2926 1338 2930 1342
rect 2966 1338 2970 1342
rect 3006 1338 3010 1342
rect 2822 1328 2826 1332
rect 2838 1328 2842 1332
rect 2958 1328 2962 1332
rect 2854 1318 2858 1322
rect 2942 1318 2946 1322
rect 2990 1318 2994 1322
rect 2758 1278 2762 1282
rect 2782 1268 2786 1272
rect 2742 1258 2746 1262
rect 2718 1248 2722 1252
rect 2766 1248 2770 1252
rect 2710 1188 2714 1192
rect 2718 1168 2722 1172
rect 2702 1148 2706 1152
rect 2750 1238 2754 1242
rect 2830 1298 2834 1302
rect 2846 1298 2850 1302
rect 3014 1298 3018 1302
rect 2918 1278 2922 1282
rect 2966 1278 2970 1282
rect 2846 1268 2850 1272
rect 2830 1248 2834 1252
rect 2814 1228 2818 1232
rect 2798 1218 2802 1222
rect 2782 1178 2786 1182
rect 2790 1168 2794 1172
rect 2662 1138 2666 1142
rect 2678 1138 2682 1142
rect 2694 1138 2698 1142
rect 2710 1138 2714 1142
rect 2742 1138 2746 1142
rect 2750 1138 2754 1142
rect 2854 1258 2858 1262
rect 2894 1268 2898 1272
rect 2998 1268 3002 1272
rect 3006 1268 3010 1272
rect 2902 1258 2906 1262
rect 2918 1258 2922 1262
rect 2942 1258 2946 1262
rect 2974 1258 2978 1262
rect 3014 1258 3018 1262
rect 2886 1248 2890 1252
rect 2814 1158 2818 1162
rect 2806 1148 2810 1152
rect 2958 1248 2962 1252
rect 2926 1238 2930 1242
rect 2966 1238 2970 1242
rect 2918 1218 2922 1222
rect 2942 1198 2946 1202
rect 3054 1428 3058 1432
rect 3030 1368 3034 1372
rect 3190 1628 3194 1632
rect 3190 1608 3194 1612
rect 3182 1588 3186 1592
rect 3118 1568 3122 1572
rect 3142 1568 3146 1572
rect 3150 1568 3154 1572
rect 3174 1568 3178 1572
rect 3166 1558 3170 1562
rect 3126 1548 3130 1552
rect 3230 1608 3234 1612
rect 3278 1558 3282 1562
rect 3302 1718 3306 1722
rect 3326 1688 3330 1692
rect 3310 1678 3314 1682
rect 3342 1678 3346 1682
rect 3294 1668 3298 1672
rect 3318 1648 3322 1652
rect 3342 1648 3346 1652
rect 3382 1688 3386 1692
rect 3358 1678 3362 1682
rect 3374 1668 3378 1672
rect 3366 1658 3370 1662
rect 3374 1658 3378 1662
rect 3358 1638 3362 1642
rect 3422 1738 3426 1742
rect 3414 1698 3418 1702
rect 3502 1808 3506 1812
rect 3494 1798 3498 1802
rect 3478 1788 3482 1792
rect 3470 1718 3474 1722
rect 3454 1688 3458 1692
rect 3430 1678 3434 1682
rect 3438 1678 3442 1682
rect 3414 1668 3418 1672
rect 3398 1658 3402 1662
rect 3430 1658 3434 1662
rect 3398 1648 3402 1652
rect 3382 1638 3386 1642
rect 3406 1638 3410 1642
rect 3350 1588 3354 1592
rect 3334 1568 3338 1572
rect 3366 1558 3370 1562
rect 3398 1558 3402 1562
rect 3230 1548 3234 1552
rect 3358 1548 3362 1552
rect 3414 1548 3418 1552
rect 3134 1538 3138 1542
rect 3102 1528 3106 1532
rect 3110 1459 3114 1463
rect 3150 1528 3154 1532
rect 3222 1538 3226 1542
rect 3214 1528 3218 1532
rect 3230 1518 3234 1522
rect 3206 1508 3210 1512
rect 3166 1488 3170 1492
rect 3166 1478 3170 1482
rect 3342 1538 3346 1542
rect 3334 1518 3338 1522
rect 3270 1508 3274 1512
rect 3302 1508 3306 1512
rect 3278 1478 3282 1482
rect 3286 1478 3290 1482
rect 3230 1468 3234 1472
rect 3182 1458 3186 1462
rect 3222 1458 3226 1462
rect 3238 1458 3242 1462
rect 3254 1458 3258 1462
rect 3262 1458 3266 1462
rect 3294 1458 3298 1462
rect 3166 1448 3170 1452
rect 3230 1448 3234 1452
rect 3150 1438 3154 1442
rect 3190 1438 3194 1442
rect 3102 1398 3106 1402
rect 3086 1358 3090 1362
rect 3166 1348 3170 1352
rect 3078 1338 3082 1342
rect 3086 1338 3090 1342
rect 3110 1338 3114 1342
rect 3070 1328 3074 1332
rect 3174 1328 3178 1332
rect 3042 1303 3046 1307
rect 3049 1303 3053 1307
rect 3086 1298 3090 1302
rect 3038 1268 3042 1272
rect 3110 1268 3114 1272
rect 3150 1268 3154 1272
rect 3166 1268 3170 1272
rect 3054 1258 3058 1262
rect 3118 1258 3122 1262
rect 3150 1238 3154 1242
rect 3126 1228 3130 1232
rect 3022 1208 3026 1212
rect 3070 1208 3074 1212
rect 3014 1198 3018 1202
rect 3270 1438 3274 1442
rect 3318 1438 3322 1442
rect 3246 1428 3250 1432
rect 3486 1708 3490 1712
rect 3534 1748 3538 1752
rect 3526 1738 3530 1742
rect 3510 1728 3514 1732
rect 3558 1728 3562 1732
rect 3518 1718 3522 1722
rect 3558 1718 3562 1722
rect 3486 1698 3490 1702
rect 3470 1668 3474 1672
rect 3454 1658 3458 1662
rect 3446 1648 3450 1652
rect 3542 1708 3546 1712
rect 3526 1698 3530 1702
rect 3502 1688 3506 1692
rect 3526 1678 3530 1682
rect 3494 1648 3498 1652
rect 3486 1628 3490 1632
rect 3494 1618 3498 1622
rect 3478 1568 3482 1572
rect 3478 1558 3482 1562
rect 3350 1518 3354 1522
rect 3422 1518 3426 1522
rect 3382 1508 3386 1512
rect 3398 1498 3402 1502
rect 3374 1478 3378 1482
rect 3398 1478 3402 1482
rect 3438 1538 3442 1542
rect 3462 1538 3466 1542
rect 3478 1528 3482 1532
rect 3446 1498 3450 1502
rect 3470 1508 3474 1512
rect 3438 1478 3442 1482
rect 3398 1468 3402 1472
rect 3414 1468 3418 1472
rect 3350 1438 3354 1442
rect 3454 1478 3458 1482
rect 3414 1448 3418 1452
rect 3366 1428 3370 1432
rect 3430 1438 3434 1442
rect 3342 1418 3346 1422
rect 3342 1398 3346 1402
rect 3206 1388 3210 1392
rect 3334 1388 3338 1392
rect 3270 1368 3274 1372
rect 3286 1358 3290 1362
rect 3230 1348 3234 1352
rect 3238 1338 3242 1342
rect 3198 1318 3202 1322
rect 3206 1318 3210 1322
rect 3214 1318 3218 1322
rect 3190 1308 3194 1312
rect 3190 1278 3194 1282
rect 3278 1338 3282 1342
rect 3246 1328 3250 1332
rect 3310 1328 3314 1332
rect 3254 1298 3258 1302
rect 3254 1288 3258 1292
rect 3270 1288 3274 1292
rect 3182 1258 3186 1262
rect 3246 1258 3250 1262
rect 3278 1258 3282 1262
rect 3190 1248 3194 1252
rect 3198 1248 3202 1252
rect 2870 1188 2874 1192
rect 3062 1188 3066 1192
rect 3158 1188 3162 1192
rect 3022 1158 3026 1162
rect 2862 1148 2866 1152
rect 2662 1128 2666 1132
rect 2654 1078 2658 1082
rect 2694 1118 2698 1122
rect 2718 1128 2722 1132
rect 2758 1128 2762 1132
rect 2774 1128 2778 1132
rect 2822 1128 2826 1132
rect 2734 1098 2738 1102
rect 2686 1078 2690 1082
rect 2702 1078 2706 1082
rect 2718 1078 2722 1082
rect 2798 1108 2802 1112
rect 2614 1068 2618 1072
rect 2686 1068 2690 1072
rect 2590 1038 2594 1042
rect 2614 978 2618 982
rect 2542 948 2546 952
rect 2598 948 2602 952
rect 2438 938 2442 942
rect 2462 938 2466 942
rect 2430 888 2434 892
rect 2510 918 2514 922
rect 2462 888 2466 892
rect 2446 878 2450 882
rect 2454 878 2458 882
rect 2470 878 2474 882
rect 2518 878 2522 882
rect 2502 868 2506 872
rect 2438 858 2442 862
rect 2494 858 2498 862
rect 2486 848 2490 852
rect 2502 848 2506 852
rect 2518 848 2522 852
rect 2470 838 2474 842
rect 2622 888 2626 892
rect 2606 868 2610 872
rect 2614 868 2618 872
rect 2582 858 2586 862
rect 2590 838 2594 842
rect 2550 818 2554 822
rect 2538 803 2542 807
rect 2545 803 2549 807
rect 2406 788 2410 792
rect 2422 788 2426 792
rect 2486 788 2490 792
rect 2414 758 2418 762
rect 2430 758 2434 762
rect 2446 758 2450 762
rect 2534 758 2538 762
rect 2406 748 2410 752
rect 2438 748 2442 752
rect 2470 748 2474 752
rect 2502 748 2506 752
rect 2550 748 2554 752
rect 2462 738 2466 742
rect 2422 728 2426 732
rect 2454 728 2458 732
rect 2494 728 2498 732
rect 2398 718 2402 722
rect 2606 788 2610 792
rect 2566 748 2570 752
rect 2374 708 2378 712
rect 2542 708 2546 712
rect 2558 708 2562 712
rect 2366 698 2370 702
rect 2326 688 2330 692
rect 2350 688 2354 692
rect 2494 688 2498 692
rect 2334 678 2338 682
rect 2398 678 2402 682
rect 2414 678 2418 682
rect 2438 678 2442 682
rect 2286 668 2290 672
rect 2366 668 2370 672
rect 2326 648 2330 652
rect 2366 648 2370 652
rect 2286 638 2290 642
rect 2318 578 2322 582
rect 2286 568 2290 572
rect 2278 558 2282 562
rect 2406 668 2410 672
rect 2390 648 2394 652
rect 2382 638 2386 642
rect 2406 638 2410 642
rect 2374 608 2378 612
rect 2374 578 2378 582
rect 2342 558 2346 562
rect 2310 548 2314 552
rect 2366 548 2370 552
rect 2302 538 2306 542
rect 2358 538 2362 542
rect 2310 528 2314 532
rect 2270 498 2274 502
rect 2142 488 2146 492
rect 2174 478 2178 482
rect 2254 478 2258 482
rect 2134 468 2138 472
rect 2182 468 2186 472
rect 2230 458 2234 462
rect 2118 408 2122 412
rect 2110 398 2114 402
rect 2166 448 2170 452
rect 2150 438 2154 442
rect 2166 428 2170 432
rect 2174 428 2178 432
rect 2142 418 2146 422
rect 2102 378 2106 382
rect 2102 338 2106 342
rect 2078 328 2082 332
rect 2118 328 2122 332
rect 2142 348 2146 352
rect 2094 278 2098 282
rect 2094 268 2098 272
rect 2110 268 2114 272
rect 2022 258 2026 262
rect 2062 258 2066 262
rect 2046 248 2050 252
rect 2062 248 2066 252
rect 2030 228 2034 232
rect 2086 258 2090 262
rect 2246 468 2250 472
rect 2302 478 2306 482
rect 2318 478 2322 482
rect 2334 478 2338 482
rect 2382 548 2386 552
rect 2390 508 2394 512
rect 2478 658 2482 662
rect 2462 648 2466 652
rect 2470 638 2474 642
rect 2510 638 2514 642
rect 2558 648 2562 652
rect 2478 618 2482 622
rect 2542 618 2546 622
rect 2430 578 2434 582
rect 2446 558 2450 562
rect 2454 548 2458 552
rect 2430 528 2434 532
rect 2350 478 2354 482
rect 2398 478 2402 482
rect 2538 603 2542 607
rect 2545 603 2549 607
rect 2558 598 2562 602
rect 2662 1058 2666 1062
rect 2686 1058 2690 1062
rect 2638 988 2642 992
rect 2806 1098 2810 1102
rect 2806 1068 2810 1072
rect 2710 1048 2714 1052
rect 2734 1048 2738 1052
rect 2742 1038 2746 1042
rect 2702 1008 2706 1012
rect 2718 1008 2722 1012
rect 2766 1058 2770 1062
rect 2782 1058 2786 1062
rect 2782 1038 2786 1042
rect 2798 1038 2802 1042
rect 2830 1108 2834 1112
rect 2838 1078 2842 1082
rect 2846 1078 2850 1082
rect 2846 1048 2850 1052
rect 2886 1138 2890 1142
rect 2902 1128 2906 1132
rect 2878 1118 2882 1122
rect 2894 1108 2898 1112
rect 2902 1098 2906 1102
rect 2894 1068 2898 1072
rect 2910 1068 2914 1072
rect 2878 1058 2882 1062
rect 2934 1138 2938 1142
rect 2926 1078 2930 1082
rect 2966 1138 2970 1142
rect 2950 1128 2954 1132
rect 2998 1138 3002 1142
rect 2998 1128 3002 1132
rect 2998 1108 3002 1112
rect 2934 1068 2938 1072
rect 2942 1058 2946 1062
rect 2958 1058 2962 1062
rect 2870 1048 2874 1052
rect 2806 1028 2810 1032
rect 2814 1028 2818 1032
rect 2822 1008 2826 1012
rect 2846 1008 2850 1012
rect 2750 978 2754 982
rect 2774 958 2778 962
rect 2806 958 2810 962
rect 2662 948 2666 952
rect 2726 948 2730 952
rect 2782 948 2786 952
rect 2774 938 2778 942
rect 2710 928 2714 932
rect 2742 928 2746 932
rect 2710 908 2714 912
rect 2742 908 2746 912
rect 2774 908 2778 912
rect 2694 898 2698 902
rect 2758 888 2762 892
rect 2742 878 2746 882
rect 2750 878 2754 882
rect 2678 868 2682 872
rect 2678 858 2682 862
rect 2654 848 2658 852
rect 2678 848 2682 852
rect 2646 818 2650 822
rect 2694 838 2698 842
rect 2710 818 2714 822
rect 2750 818 2754 822
rect 2678 808 2682 812
rect 2646 778 2650 782
rect 2630 768 2634 772
rect 2742 768 2746 772
rect 2638 758 2642 762
rect 2622 748 2626 752
rect 2614 738 2618 742
rect 2622 738 2626 742
rect 2606 728 2610 732
rect 2630 728 2634 732
rect 2614 718 2618 722
rect 2710 748 2714 752
rect 2654 738 2658 742
rect 2662 728 2666 732
rect 2726 728 2730 732
rect 2654 688 2658 692
rect 2662 688 2666 692
rect 2710 688 2714 692
rect 2742 738 2746 742
rect 2742 718 2746 722
rect 2734 708 2738 712
rect 2766 878 2770 882
rect 2798 918 2802 922
rect 2830 998 2834 1002
rect 2854 958 2858 962
rect 2830 938 2834 942
rect 2846 928 2850 932
rect 2814 888 2818 892
rect 2822 888 2826 892
rect 2902 1048 2906 1052
rect 2902 968 2906 972
rect 2942 1048 2946 1052
rect 2942 1028 2946 1032
rect 3014 1128 3018 1132
rect 3006 1098 3010 1102
rect 2998 1068 3002 1072
rect 2990 1058 2994 1062
rect 2942 1008 2946 1012
rect 2950 1008 2954 1012
rect 2974 1008 2978 1012
rect 3042 1103 3046 1107
rect 3049 1103 3053 1107
rect 3030 1098 3034 1102
rect 3086 1168 3090 1172
rect 3110 1148 3114 1152
rect 3150 1148 3154 1152
rect 3062 1048 3066 1052
rect 3022 1028 3026 1032
rect 3046 1028 3050 1032
rect 3014 998 3018 1002
rect 3046 988 3050 992
rect 2918 978 2922 982
rect 2942 978 2946 982
rect 2894 938 2898 942
rect 2958 958 2962 962
rect 2926 948 2930 952
rect 2934 948 2938 952
rect 2974 948 2978 952
rect 2998 948 3002 952
rect 2982 938 2986 942
rect 3054 938 3058 942
rect 2918 928 2922 932
rect 2950 928 2954 932
rect 2966 928 2970 932
rect 2862 908 2866 912
rect 2878 908 2882 912
rect 2790 878 2794 882
rect 2798 878 2802 882
rect 2854 878 2858 882
rect 2958 898 2962 902
rect 2982 908 2986 912
rect 2974 898 2978 902
rect 2942 888 2946 892
rect 2902 878 2906 882
rect 2926 878 2930 882
rect 2782 858 2786 862
rect 2838 858 2842 862
rect 2862 858 2866 862
rect 2926 858 2930 862
rect 2934 858 2938 862
rect 2774 838 2778 842
rect 2878 848 2882 852
rect 2910 848 2914 852
rect 2806 818 2810 822
rect 2830 818 2834 822
rect 2782 798 2786 802
rect 2798 788 2802 792
rect 2782 768 2786 772
rect 2766 748 2770 752
rect 2774 748 2778 752
rect 2790 738 2794 742
rect 2758 688 2762 692
rect 2622 678 2626 682
rect 2694 678 2698 682
rect 2726 678 2730 682
rect 2742 678 2746 682
rect 2646 668 2650 672
rect 2678 668 2682 672
rect 2766 668 2770 672
rect 2630 638 2634 642
rect 2686 648 2690 652
rect 2702 648 2706 652
rect 2742 648 2746 652
rect 2934 838 2938 842
rect 2886 818 2890 822
rect 3042 903 3046 907
rect 3049 903 3053 907
rect 2990 888 2994 892
rect 3038 888 3042 892
rect 3030 878 3034 882
rect 3054 878 3058 882
rect 2990 848 2994 852
rect 2950 808 2954 812
rect 2854 778 2858 782
rect 2958 778 2962 782
rect 2966 778 2970 782
rect 2846 748 2850 752
rect 2894 747 2898 751
rect 2822 728 2826 732
rect 2790 718 2794 722
rect 2806 718 2810 722
rect 2774 638 2778 642
rect 2670 618 2674 622
rect 2622 608 2626 612
rect 2558 578 2562 582
rect 2654 578 2658 582
rect 2582 558 2586 562
rect 2598 558 2602 562
rect 2646 558 2650 562
rect 2686 558 2690 562
rect 2734 558 2738 562
rect 2510 548 2514 552
rect 2502 538 2506 542
rect 2542 538 2546 542
rect 2582 538 2586 542
rect 2494 518 2498 522
rect 2486 508 2490 512
rect 2566 528 2570 532
rect 2510 498 2514 502
rect 2350 468 2354 472
rect 2430 468 2434 472
rect 2294 458 2298 462
rect 2310 458 2314 462
rect 2318 458 2322 462
rect 2238 448 2242 452
rect 2246 448 2250 452
rect 2302 448 2306 452
rect 2246 408 2250 412
rect 2230 398 2234 402
rect 2206 378 2210 382
rect 2318 438 2322 442
rect 2302 428 2306 432
rect 2182 358 2186 362
rect 2206 358 2210 362
rect 2254 358 2258 362
rect 2278 358 2282 362
rect 2342 458 2346 462
rect 2350 458 2354 462
rect 2334 448 2338 452
rect 2374 438 2378 442
rect 2326 408 2330 412
rect 2350 408 2354 412
rect 2366 408 2370 412
rect 2366 398 2370 402
rect 2358 378 2362 382
rect 2198 348 2202 352
rect 2238 348 2242 352
rect 2174 338 2178 342
rect 2206 338 2210 342
rect 2190 328 2194 332
rect 2158 308 2162 312
rect 2262 328 2266 332
rect 2302 338 2306 342
rect 2310 328 2314 332
rect 2326 328 2330 332
rect 2222 318 2226 322
rect 2278 318 2282 322
rect 2254 308 2258 312
rect 2150 298 2154 302
rect 2166 298 2170 302
rect 2454 458 2458 462
rect 2390 418 2394 422
rect 2430 438 2434 442
rect 2502 448 2506 452
rect 2454 428 2458 432
rect 2446 418 2450 422
rect 2470 398 2474 402
rect 2454 378 2458 382
rect 2430 358 2434 362
rect 2382 348 2386 352
rect 2342 298 2346 302
rect 2286 288 2290 292
rect 2198 278 2202 282
rect 2294 278 2298 282
rect 2134 268 2138 272
rect 2214 268 2218 272
rect 2302 268 2306 272
rect 2318 268 2322 272
rect 2326 268 2330 272
rect 2150 258 2154 262
rect 2222 258 2226 262
rect 2254 258 2258 262
rect 2078 218 2082 222
rect 2054 158 2058 162
rect 2078 158 2082 162
rect 2046 148 2050 152
rect 1910 138 1914 142
rect 1886 128 1890 132
rect 1934 128 1938 132
rect 1926 118 1930 122
rect 1846 78 1850 82
rect 1870 78 1874 82
rect 1886 78 1890 82
rect 1894 78 1898 82
rect 1942 108 1946 112
rect 1942 98 1946 102
rect 1918 78 1922 82
rect 2094 248 2098 252
rect 2110 248 2114 252
rect 2238 248 2242 252
rect 2270 248 2274 252
rect 2286 248 2290 252
rect 2206 238 2210 242
rect 2254 238 2258 242
rect 2126 228 2130 232
rect 2158 228 2162 232
rect 2126 158 2130 162
rect 2166 178 2170 182
rect 2318 228 2322 232
rect 2334 228 2338 232
rect 2286 218 2290 222
rect 2294 218 2298 222
rect 2278 198 2282 202
rect 2254 158 2258 162
rect 2110 148 2114 152
rect 2142 148 2146 152
rect 2166 148 2170 152
rect 2190 148 2194 152
rect 2206 148 2210 152
rect 2398 338 2402 342
rect 2430 348 2434 352
rect 2446 348 2450 352
rect 2422 338 2426 342
rect 2438 338 2442 342
rect 2414 328 2418 332
rect 2374 308 2378 312
rect 2502 418 2506 422
rect 2526 518 2530 522
rect 2558 488 2562 492
rect 2566 478 2570 482
rect 2534 448 2538 452
rect 2478 368 2482 372
rect 2538 403 2542 407
rect 2545 403 2549 407
rect 2550 358 2554 362
rect 2510 338 2514 342
rect 2462 328 2466 332
rect 2494 328 2498 332
rect 2486 318 2490 322
rect 2470 308 2474 312
rect 2422 298 2426 302
rect 2502 298 2506 302
rect 2534 338 2538 342
rect 2358 288 2362 292
rect 2518 288 2522 292
rect 2430 278 2434 282
rect 2542 298 2546 302
rect 2406 268 2410 272
rect 2470 268 2474 272
rect 2494 268 2498 272
rect 2510 268 2514 272
rect 2518 268 2522 272
rect 2382 258 2386 262
rect 2446 258 2450 262
rect 2398 248 2402 252
rect 2430 248 2434 252
rect 2478 248 2482 252
rect 2398 238 2402 242
rect 2470 238 2474 242
rect 2350 208 2354 212
rect 2342 178 2346 182
rect 2382 208 2386 212
rect 2390 208 2394 212
rect 2382 178 2386 182
rect 2302 158 2306 162
rect 2350 158 2354 162
rect 2294 148 2298 152
rect 2326 148 2330 152
rect 2358 148 2362 152
rect 2078 138 2082 142
rect 2118 138 2122 142
rect 2158 138 2162 142
rect 2206 138 2210 142
rect 2230 138 2234 142
rect 2270 138 2274 142
rect 1974 118 1978 122
rect 1974 98 1978 102
rect 1958 78 1962 82
rect 1982 78 1986 82
rect 2006 118 2010 122
rect 2026 103 2030 107
rect 2033 103 2037 107
rect 2046 98 2050 102
rect 2014 78 2018 82
rect 2030 78 2034 82
rect 2046 78 2050 82
rect 2070 128 2074 132
rect 2110 128 2114 132
rect 2142 128 2146 132
rect 2150 128 2154 132
rect 2166 128 2170 132
rect 2110 118 2114 122
rect 2182 118 2186 122
rect 2094 108 2098 112
rect 2062 78 2066 82
rect 2190 108 2194 112
rect 2254 108 2258 112
rect 2286 98 2290 102
rect 2294 98 2298 102
rect 2510 218 2514 222
rect 2542 258 2546 262
rect 2558 328 2562 332
rect 2606 528 2610 532
rect 2590 508 2594 512
rect 2622 538 2626 542
rect 2614 508 2618 512
rect 2630 528 2634 532
rect 2678 548 2682 552
rect 2718 548 2722 552
rect 2686 538 2690 542
rect 2654 518 2658 522
rect 2678 518 2682 522
rect 2662 498 2666 502
rect 2654 488 2658 492
rect 2662 488 2666 492
rect 2646 478 2650 482
rect 2606 468 2610 472
rect 2670 468 2674 472
rect 2590 428 2594 432
rect 2574 398 2578 402
rect 2582 348 2586 352
rect 2606 368 2610 372
rect 2758 558 2762 562
rect 2774 558 2778 562
rect 2742 548 2746 552
rect 2742 538 2746 542
rect 2702 528 2706 532
rect 2726 528 2730 532
rect 2702 518 2706 522
rect 2694 508 2698 512
rect 2774 498 2778 502
rect 2806 708 2810 712
rect 2814 698 2818 702
rect 2958 738 2962 742
rect 2854 728 2858 732
rect 2862 718 2866 722
rect 2854 698 2858 702
rect 2798 658 2802 662
rect 2814 658 2818 662
rect 2838 658 2842 662
rect 2846 638 2850 642
rect 2974 748 2978 752
rect 2894 708 2898 712
rect 2958 708 2962 712
rect 2982 708 2986 712
rect 2870 678 2874 682
rect 2998 838 3002 842
rect 3014 838 3018 842
rect 3094 1138 3098 1142
rect 3134 1138 3138 1142
rect 3150 1138 3154 1142
rect 3110 1128 3114 1132
rect 3174 1168 3178 1172
rect 3174 1148 3178 1152
rect 3190 1148 3194 1152
rect 3214 1138 3218 1142
rect 3182 1128 3186 1132
rect 3198 1128 3202 1132
rect 3214 1128 3218 1132
rect 3230 1128 3234 1132
rect 3238 1128 3242 1132
rect 3166 1118 3170 1122
rect 3238 1118 3242 1122
rect 3262 1118 3266 1122
rect 3158 1108 3162 1112
rect 3214 1108 3218 1112
rect 3126 1098 3130 1102
rect 3086 1088 3090 1092
rect 3118 1078 3122 1082
rect 3150 1078 3154 1082
rect 3158 1078 3162 1082
rect 3206 1078 3210 1082
rect 3102 1058 3106 1062
rect 3086 1038 3090 1042
rect 3078 1018 3082 1022
rect 3110 978 3114 982
rect 3070 948 3074 952
rect 3102 948 3106 952
rect 3078 938 3082 942
rect 3078 928 3082 932
rect 3166 1068 3170 1072
rect 3174 1068 3178 1072
rect 3126 1058 3130 1062
rect 3150 1048 3154 1052
rect 3246 1068 3250 1072
rect 3230 1058 3234 1062
rect 3198 1048 3202 1052
rect 3254 1048 3258 1052
rect 3182 1038 3186 1042
rect 3198 1038 3202 1042
rect 3142 1018 3146 1022
rect 3182 1008 3186 1012
rect 3134 988 3138 992
rect 3166 988 3170 992
rect 3150 958 3154 962
rect 3142 948 3146 952
rect 3174 938 3178 942
rect 3126 928 3130 932
rect 3102 918 3106 922
rect 3118 918 3122 922
rect 3078 878 3082 882
rect 3102 878 3106 882
rect 3062 828 3066 832
rect 3166 928 3170 932
rect 3166 918 3170 922
rect 3206 1028 3210 1032
rect 3230 1028 3234 1032
rect 3262 1028 3266 1032
rect 3198 998 3202 1002
rect 3190 958 3194 962
rect 3286 1248 3290 1252
rect 3294 1218 3298 1222
rect 3382 1418 3386 1422
rect 3350 1338 3354 1342
rect 3350 1328 3354 1332
rect 3406 1388 3410 1392
rect 3374 1328 3378 1332
rect 3406 1328 3410 1332
rect 3366 1298 3370 1302
rect 3374 1298 3378 1302
rect 3454 1418 3458 1422
rect 3438 1338 3442 1342
rect 3518 1628 3522 1632
rect 3510 1598 3514 1602
rect 3510 1588 3514 1592
rect 3510 1568 3514 1572
rect 3494 1528 3498 1532
rect 3502 1528 3506 1532
rect 3526 1608 3530 1612
rect 3550 1558 3554 1562
rect 3542 1548 3546 1552
rect 3486 1488 3490 1492
rect 3502 1478 3506 1482
rect 3542 1478 3546 1482
rect 3518 1468 3522 1472
rect 3494 1458 3498 1462
rect 3470 1448 3474 1452
rect 3454 1408 3458 1412
rect 3462 1408 3466 1412
rect 3558 1448 3562 1452
rect 3550 1438 3554 1442
rect 3542 1418 3546 1422
rect 3542 1408 3546 1412
rect 3470 1378 3474 1382
rect 3534 1378 3538 1382
rect 3502 1368 3506 1372
rect 3526 1368 3530 1372
rect 3478 1358 3482 1362
rect 3510 1358 3514 1362
rect 3454 1338 3458 1342
rect 3470 1338 3474 1342
rect 3494 1338 3498 1342
rect 3534 1338 3538 1342
rect 3542 1338 3546 1342
rect 3470 1328 3474 1332
rect 3486 1328 3490 1332
rect 3462 1318 3466 1322
rect 3446 1308 3450 1312
rect 3478 1288 3482 1292
rect 3374 1278 3378 1282
rect 3406 1278 3410 1282
rect 3414 1278 3418 1282
rect 3310 1258 3314 1262
rect 3342 1258 3346 1262
rect 3358 1258 3362 1262
rect 3398 1258 3402 1262
rect 3350 1248 3354 1252
rect 3374 1248 3378 1252
rect 3390 1248 3394 1252
rect 3342 1228 3346 1232
rect 3326 1218 3330 1222
rect 3302 1168 3306 1172
rect 3422 1268 3426 1272
rect 3446 1268 3450 1272
rect 3558 1268 3562 1272
rect 3430 1258 3434 1262
rect 3398 1178 3402 1182
rect 3446 1168 3450 1172
rect 3342 1148 3346 1152
rect 3366 1158 3370 1162
rect 3374 1158 3378 1162
rect 3406 1158 3410 1162
rect 3462 1158 3466 1162
rect 3326 1138 3330 1142
rect 3342 1138 3346 1142
rect 3382 1138 3386 1142
rect 3278 1108 3282 1112
rect 3294 1098 3298 1102
rect 3286 1088 3290 1092
rect 3310 1098 3314 1102
rect 3382 1088 3386 1092
rect 3334 1078 3338 1082
rect 3286 1058 3290 1062
rect 3326 1058 3330 1062
rect 3334 1048 3338 1052
rect 3430 1148 3434 1152
rect 3494 1248 3498 1252
rect 3558 1168 3562 1172
rect 3526 1148 3530 1152
rect 3430 1088 3434 1092
rect 3494 1098 3498 1102
rect 3406 1058 3410 1062
rect 3358 1048 3362 1052
rect 3366 1048 3370 1052
rect 3398 1048 3402 1052
rect 3462 1048 3466 1052
rect 3318 1038 3322 1042
rect 3350 1038 3354 1042
rect 3406 1038 3410 1042
rect 3270 1008 3274 1012
rect 3302 968 3306 972
rect 3350 968 3354 972
rect 3206 948 3210 952
rect 3230 948 3234 952
rect 3238 948 3242 952
rect 3190 938 3194 942
rect 3214 938 3218 942
rect 3246 938 3250 942
rect 3278 938 3282 942
rect 3246 928 3250 932
rect 3254 908 3258 912
rect 3342 958 3346 962
rect 3310 938 3314 942
rect 3350 928 3354 932
rect 3414 1008 3418 1012
rect 3390 968 3394 972
rect 3406 968 3410 972
rect 3382 948 3386 952
rect 3390 948 3394 952
rect 3374 928 3378 932
rect 3406 928 3410 932
rect 3382 918 3386 922
rect 3406 918 3410 922
rect 3390 908 3394 912
rect 3206 888 3210 892
rect 3342 888 3346 892
rect 3166 878 3170 882
rect 3222 878 3226 882
rect 3278 878 3282 882
rect 3334 878 3338 882
rect 3390 878 3394 882
rect 3286 858 3290 862
rect 3342 858 3346 862
rect 3086 848 3090 852
rect 3126 848 3130 852
rect 3134 848 3138 852
rect 3174 848 3178 852
rect 3230 848 3234 852
rect 3126 838 3130 842
rect 3078 808 3082 812
rect 3254 818 3258 822
rect 3422 988 3426 992
rect 3462 958 3466 962
rect 3430 948 3434 952
rect 3446 938 3450 942
rect 3406 858 3410 862
rect 3414 858 3418 862
rect 3134 798 3138 802
rect 3374 798 3378 802
rect 3398 798 3402 802
rect 3214 778 3218 782
rect 3086 768 3090 772
rect 3102 768 3106 772
rect 3142 768 3146 772
rect 3102 758 3106 762
rect 3038 748 3042 752
rect 3062 748 3066 752
rect 3006 738 3010 742
rect 3030 738 3034 742
rect 3054 728 3058 732
rect 2998 708 3002 712
rect 2990 698 2994 702
rect 3030 708 3034 712
rect 2926 688 2930 692
rect 3014 688 3018 692
rect 3006 678 3010 682
rect 3022 678 3026 682
rect 2878 668 2882 672
rect 2950 668 2954 672
rect 2974 668 2978 672
rect 2862 588 2866 592
rect 2862 578 2866 582
rect 2894 658 2898 662
rect 2902 658 2906 662
rect 2926 648 2930 652
rect 2886 638 2890 642
rect 2902 638 2906 642
rect 2870 568 2874 572
rect 2806 548 2810 552
rect 2806 538 2810 542
rect 2806 518 2810 522
rect 2814 498 2818 502
rect 2838 498 2842 502
rect 2710 488 2714 492
rect 2734 488 2738 492
rect 2774 488 2778 492
rect 2790 488 2794 492
rect 2814 488 2818 492
rect 2718 478 2722 482
rect 2742 478 2746 482
rect 2766 478 2770 482
rect 2790 478 2794 482
rect 2806 478 2810 482
rect 2638 458 2642 462
rect 2654 448 2658 452
rect 2686 448 2690 452
rect 2622 418 2626 422
rect 2614 358 2618 362
rect 2750 448 2754 452
rect 2718 438 2722 442
rect 2750 438 2754 442
rect 2758 438 2762 442
rect 2678 368 2682 372
rect 2678 358 2682 362
rect 2622 348 2626 352
rect 2654 348 2658 352
rect 2574 338 2578 342
rect 2622 338 2626 342
rect 2638 338 2642 342
rect 2686 338 2690 342
rect 2574 318 2578 322
rect 2590 298 2594 302
rect 2558 238 2562 242
rect 2550 218 2554 222
rect 2538 203 2542 207
rect 2545 203 2549 207
rect 2590 248 2594 252
rect 2590 238 2594 242
rect 2526 198 2530 202
rect 2566 198 2570 202
rect 2438 158 2442 162
rect 2446 158 2450 162
rect 2422 148 2426 152
rect 2502 148 2506 152
rect 2630 298 2634 302
rect 2638 278 2642 282
rect 2622 268 2626 272
rect 2630 268 2634 272
rect 2670 268 2674 272
rect 2614 238 2618 242
rect 2606 178 2610 182
rect 2422 138 2426 142
rect 2438 138 2442 142
rect 2486 138 2490 142
rect 2510 138 2514 142
rect 2406 128 2410 132
rect 2422 128 2426 132
rect 2334 108 2338 112
rect 2350 108 2354 112
rect 2374 108 2378 112
rect 2398 98 2402 102
rect 2414 98 2418 102
rect 2126 88 2130 92
rect 2190 78 2194 82
rect 2158 68 2162 72
rect 2206 68 2210 72
rect 2230 68 2234 72
rect 2262 68 2266 72
rect 2286 68 2290 72
rect 1998 58 2002 62
rect 2118 58 2122 62
rect 2142 58 2146 62
rect 1838 48 1842 52
rect 1910 48 1914 52
rect 1950 48 1954 52
rect 1830 38 1834 42
rect 1846 38 1850 42
rect 1870 38 1874 42
rect 1990 38 1994 42
rect 2214 58 2218 62
rect 2238 58 2242 62
rect 2254 58 2258 62
rect 2206 18 2210 22
rect 2318 68 2322 72
rect 2326 58 2330 62
rect 2366 58 2370 62
rect 2390 58 2394 62
rect 2334 48 2338 52
rect 2374 48 2378 52
rect 2406 48 2410 52
rect 2302 38 2306 42
rect 2358 28 2362 32
rect 2494 128 2498 132
rect 2478 118 2482 122
rect 2446 98 2450 102
rect 2454 98 2458 102
rect 2566 118 2570 122
rect 2662 258 2666 262
rect 2678 238 2682 242
rect 2718 338 2722 342
rect 2742 348 2746 352
rect 2750 318 2754 322
rect 2798 438 2802 442
rect 2830 478 2834 482
rect 2870 528 2874 532
rect 2846 458 2850 462
rect 2790 408 2794 412
rect 2814 408 2818 412
rect 2862 428 2866 432
rect 2830 398 2834 402
rect 2814 368 2818 372
rect 2782 348 2786 352
rect 2806 348 2810 352
rect 2774 338 2778 342
rect 2838 348 2842 352
rect 2926 618 2930 622
rect 2934 618 2938 622
rect 2886 538 2890 542
rect 2926 558 2930 562
rect 2910 548 2914 552
rect 2926 538 2930 542
rect 2910 528 2914 532
rect 2958 628 2962 632
rect 2990 638 2994 642
rect 2974 618 2978 622
rect 3042 703 3046 707
rect 3049 703 3053 707
rect 3038 678 3042 682
rect 3046 638 3050 642
rect 3030 618 3034 622
rect 2998 608 3002 612
rect 3022 608 3026 612
rect 2990 598 2994 602
rect 2958 568 2962 572
rect 2966 558 2970 562
rect 2998 558 3002 562
rect 2950 548 2954 552
rect 2950 528 2954 532
rect 2982 548 2986 552
rect 2998 548 3002 552
rect 3014 548 3018 552
rect 3006 538 3010 542
rect 2998 508 3002 512
rect 2934 468 2938 472
rect 2878 448 2882 452
rect 2910 458 2914 462
rect 2958 458 2962 462
rect 2990 458 2994 462
rect 2894 448 2898 452
rect 2926 448 2930 452
rect 2886 428 2890 432
rect 2870 408 2874 412
rect 2902 408 2906 412
rect 2966 418 2970 422
rect 2950 398 2954 402
rect 2950 388 2954 392
rect 2862 368 2866 372
rect 2870 348 2874 352
rect 2886 348 2890 352
rect 2958 348 2962 352
rect 2854 338 2858 342
rect 2790 318 2794 322
rect 2806 318 2810 322
rect 2822 318 2826 322
rect 2838 318 2842 322
rect 2750 308 2754 312
rect 2766 308 2770 312
rect 2734 288 2738 292
rect 2710 278 2714 282
rect 2718 268 2722 272
rect 2702 258 2706 262
rect 2894 338 2898 342
rect 2902 338 2906 342
rect 2942 338 2946 342
rect 2950 328 2954 332
rect 2958 328 2962 332
rect 2894 308 2898 312
rect 2998 408 3002 412
rect 2998 388 3002 392
rect 3006 368 3010 372
rect 2998 338 3002 342
rect 2990 328 2994 332
rect 2910 308 2914 312
rect 2918 308 2922 312
rect 2958 308 2962 312
rect 2982 308 2986 312
rect 2990 298 2994 302
rect 2878 288 2882 292
rect 2918 288 2922 292
rect 2822 278 2826 282
rect 2806 268 2810 272
rect 2846 268 2850 272
rect 2726 258 2730 262
rect 2750 258 2754 262
rect 2782 258 2786 262
rect 2806 258 2810 262
rect 2822 258 2826 262
rect 2710 238 2714 242
rect 2694 208 2698 212
rect 2718 218 2722 222
rect 2742 198 2746 202
rect 2726 188 2730 192
rect 2662 158 2666 162
rect 2710 158 2714 162
rect 2654 148 2658 152
rect 2646 128 2650 132
rect 2622 118 2626 122
rect 2654 118 2658 122
rect 2606 98 2610 102
rect 2614 98 2618 102
rect 2502 88 2506 92
rect 2566 88 2570 92
rect 2590 88 2594 92
rect 2438 78 2442 82
rect 2462 78 2466 82
rect 2478 78 2482 82
rect 2558 68 2562 72
rect 2438 58 2442 62
rect 2454 58 2458 62
rect 2462 58 2466 62
rect 2430 48 2434 52
rect 2422 18 2426 22
rect 2334 8 2338 12
rect 2366 8 2370 12
rect 2414 8 2418 12
rect 2542 58 2546 62
rect 2550 48 2554 52
rect 2590 68 2594 72
rect 2614 78 2618 82
rect 2630 78 2634 82
rect 2662 108 2666 112
rect 2646 68 2650 72
rect 2694 128 2698 132
rect 2670 98 2674 102
rect 2678 98 2682 102
rect 2718 88 2722 92
rect 2694 78 2698 82
rect 2734 158 2738 162
rect 2790 248 2794 252
rect 2774 218 2778 222
rect 2758 178 2762 182
rect 2934 278 2938 282
rect 2950 278 2954 282
rect 2974 278 2978 282
rect 2902 268 2906 272
rect 2926 268 2930 272
rect 2854 258 2858 262
rect 2870 258 2874 262
rect 2862 228 2866 232
rect 2870 228 2874 232
rect 2846 198 2850 202
rect 2838 158 2842 162
rect 2886 258 2890 262
rect 2886 228 2890 232
rect 2934 258 2938 262
rect 2950 248 2954 252
rect 2942 238 2946 242
rect 2958 208 2962 212
rect 3054 598 3058 602
rect 3262 768 3266 772
rect 3158 758 3162 762
rect 3182 758 3186 762
rect 3214 758 3218 762
rect 3190 748 3194 752
rect 3222 748 3226 752
rect 3286 748 3290 752
rect 3118 738 3122 742
rect 3198 738 3202 742
rect 3174 728 3178 732
rect 3230 728 3234 732
rect 3110 708 3114 712
rect 3142 708 3146 712
rect 3158 708 3162 712
rect 3198 718 3202 722
rect 3198 708 3202 712
rect 3206 698 3210 702
rect 3110 688 3114 692
rect 3158 688 3162 692
rect 3078 678 3082 682
rect 3094 678 3098 682
rect 3110 678 3114 682
rect 3078 668 3082 672
rect 3070 658 3074 662
rect 3062 578 3066 582
rect 3118 668 3122 672
rect 3150 668 3154 672
rect 3222 668 3226 672
rect 3110 658 3114 662
rect 3126 658 3130 662
rect 3166 658 3170 662
rect 3182 658 3186 662
rect 3206 658 3210 662
rect 3102 628 3106 632
rect 3110 598 3114 602
rect 3086 568 3090 572
rect 3110 568 3114 572
rect 3030 558 3034 562
rect 3046 558 3050 562
rect 3038 538 3042 542
rect 3042 503 3046 507
rect 3049 503 3053 507
rect 3038 478 3042 482
rect 3030 438 3034 442
rect 3030 368 3034 372
rect 3030 338 3034 342
rect 3006 288 3010 292
rect 2998 268 3002 272
rect 3006 268 3010 272
rect 2926 178 2930 182
rect 2950 168 2954 172
rect 2910 158 2914 162
rect 2918 158 2922 162
rect 2942 158 2946 162
rect 2806 148 2810 152
rect 2830 148 2834 152
rect 2854 148 2858 152
rect 2750 128 2754 132
rect 2878 148 2882 152
rect 2774 138 2778 142
rect 2886 138 2890 142
rect 2902 138 2906 142
rect 2806 128 2810 132
rect 2830 128 2834 132
rect 2766 118 2770 122
rect 2790 118 2794 122
rect 2774 108 2778 112
rect 2758 88 2762 92
rect 2678 68 2682 72
rect 2726 68 2730 72
rect 2750 68 2754 72
rect 2670 58 2674 62
rect 2702 58 2706 62
rect 2718 58 2722 62
rect 2734 58 2738 62
rect 2774 58 2778 62
rect 2894 108 2898 112
rect 2974 188 2978 192
rect 3102 558 3106 562
rect 3070 548 3074 552
rect 3086 538 3090 542
rect 3094 518 3098 522
rect 3070 488 3074 492
rect 3094 488 3098 492
rect 3110 518 3114 522
rect 3102 468 3106 472
rect 3110 468 3114 472
rect 3110 458 3114 462
rect 3086 448 3090 452
rect 3110 448 3114 452
rect 3078 438 3082 442
rect 3262 659 3266 663
rect 3326 728 3330 732
rect 3334 708 3338 712
rect 3310 688 3314 692
rect 3358 698 3362 702
rect 3366 678 3370 682
rect 3326 668 3330 672
rect 3318 658 3322 662
rect 3134 638 3138 642
rect 3190 638 3194 642
rect 3214 638 3218 642
rect 3342 618 3346 622
rect 3286 588 3290 592
rect 3142 568 3146 572
rect 3238 558 3242 562
rect 3158 548 3162 552
rect 3182 548 3186 552
rect 3198 548 3202 552
rect 3230 548 3234 552
rect 3278 548 3282 552
rect 3318 548 3322 552
rect 3190 528 3194 532
rect 3222 528 3226 532
rect 3150 498 3154 502
rect 3182 518 3186 522
rect 3198 518 3202 522
rect 3214 518 3218 522
rect 3198 508 3202 512
rect 3294 538 3298 542
rect 3326 538 3330 542
rect 3342 538 3346 542
rect 3246 528 3250 532
rect 3230 498 3234 502
rect 3278 498 3282 502
rect 3222 488 3226 492
rect 3246 478 3250 482
rect 3390 738 3394 742
rect 3422 848 3426 852
rect 3470 808 3474 812
rect 3518 1088 3522 1092
rect 3558 1048 3562 1052
rect 3526 998 3530 1002
rect 3558 998 3562 1002
rect 3526 948 3530 952
rect 3494 868 3498 872
rect 3526 868 3530 872
rect 3526 848 3530 852
rect 3558 848 3562 852
rect 3494 828 3498 832
rect 3502 788 3506 792
rect 3518 788 3522 792
rect 3558 788 3562 792
rect 3478 778 3482 782
rect 3478 758 3482 762
rect 3550 768 3554 772
rect 3438 748 3442 752
rect 3446 748 3450 752
rect 3430 728 3434 732
rect 3422 708 3426 712
rect 3422 688 3426 692
rect 3454 718 3458 722
rect 3510 688 3514 692
rect 3526 688 3530 692
rect 3414 668 3418 672
rect 3358 648 3362 652
rect 3366 638 3370 642
rect 3406 588 3410 592
rect 3422 558 3426 562
rect 3374 528 3378 532
rect 3334 478 3338 482
rect 3142 468 3146 472
rect 3206 468 3210 472
rect 3230 468 3234 472
rect 3278 468 3282 472
rect 3310 468 3314 472
rect 3334 468 3338 472
rect 3086 428 3090 432
rect 3126 428 3130 432
rect 3134 428 3138 432
rect 3142 428 3146 432
rect 3062 418 3066 422
rect 3086 418 3090 422
rect 3078 408 3082 412
rect 3086 408 3090 412
rect 3070 348 3074 352
rect 3110 368 3114 372
rect 3094 348 3098 352
rect 3118 348 3122 352
rect 3070 328 3074 332
rect 3054 318 3058 322
rect 3042 303 3046 307
rect 3049 303 3053 307
rect 3070 318 3074 322
rect 3166 448 3170 452
rect 3158 418 3162 422
rect 3150 388 3154 392
rect 3174 428 3178 432
rect 3190 418 3194 422
rect 3182 388 3186 392
rect 3158 368 3162 372
rect 3158 348 3162 352
rect 3126 338 3130 342
rect 3102 318 3106 322
rect 3142 308 3146 312
rect 3166 308 3170 312
rect 3190 368 3194 372
rect 3198 368 3202 372
rect 3262 438 3266 442
rect 3326 458 3330 462
rect 3278 448 3282 452
rect 3302 448 3306 452
rect 3286 438 3290 442
rect 3294 418 3298 422
rect 3246 388 3250 392
rect 3270 388 3274 392
rect 3246 378 3250 382
rect 3286 378 3290 382
rect 3190 348 3194 352
rect 3214 348 3218 352
rect 3198 318 3202 322
rect 3174 298 3178 302
rect 3126 278 3130 282
rect 3174 278 3178 282
rect 3238 338 3242 342
rect 3334 428 3338 432
rect 3302 388 3306 392
rect 3318 348 3322 352
rect 3366 468 3370 472
rect 3374 458 3378 462
rect 3518 658 3522 662
rect 3454 648 3458 652
rect 3526 638 3530 642
rect 3510 548 3514 552
rect 3486 538 3490 542
rect 3494 538 3498 542
rect 3390 488 3394 492
rect 3406 478 3410 482
rect 3518 528 3522 532
rect 3366 448 3370 452
rect 3342 418 3346 422
rect 3398 438 3402 442
rect 3422 418 3426 422
rect 3406 378 3410 382
rect 3382 358 3386 362
rect 3342 348 3346 352
rect 3350 338 3354 342
rect 3374 338 3378 342
rect 3398 338 3402 342
rect 3414 338 3418 342
rect 3222 328 3226 332
rect 3246 328 3250 332
rect 3262 328 3266 332
rect 3286 328 3290 332
rect 3294 328 3298 332
rect 3318 328 3322 332
rect 3254 318 3258 322
rect 3238 278 3242 282
rect 3270 298 3274 302
rect 3262 278 3266 282
rect 3142 268 3146 272
rect 3158 268 3162 272
rect 3062 248 3066 252
rect 3094 248 3098 252
rect 3078 238 3082 242
rect 3022 228 3026 232
rect 2990 188 2994 192
rect 3022 188 3026 192
rect 3046 188 3050 192
rect 3238 258 3242 262
rect 3126 248 3130 252
rect 3166 248 3170 252
rect 3150 238 3154 242
rect 3110 168 3114 172
rect 3150 168 3154 172
rect 3190 168 3194 172
rect 3062 158 3066 162
rect 3142 158 3146 162
rect 3038 148 3042 152
rect 3046 148 3050 152
rect 3094 148 3098 152
rect 2982 138 2986 142
rect 3094 138 3098 142
rect 2966 118 2970 122
rect 3006 98 3010 102
rect 3022 128 3026 132
rect 3110 128 3114 132
rect 3118 128 3122 132
rect 3042 103 3046 107
rect 3049 103 3053 107
rect 3062 98 3066 102
rect 3094 98 3098 102
rect 3014 88 3018 92
rect 3214 248 3218 252
rect 3222 228 3226 232
rect 3238 208 3242 212
rect 3230 178 3234 182
rect 3222 168 3226 172
rect 3166 158 3170 162
rect 3214 158 3218 162
rect 3174 148 3178 152
rect 3182 138 3186 142
rect 3158 118 3162 122
rect 3150 108 3154 112
rect 3174 108 3178 112
rect 3134 88 3138 92
rect 3222 118 3226 122
rect 3190 88 3194 92
rect 2806 78 2810 82
rect 2862 78 2866 82
rect 2918 78 2922 82
rect 3030 78 3034 82
rect 3046 78 3050 82
rect 2806 68 2810 72
rect 2934 68 2938 72
rect 2942 68 2946 72
rect 2950 68 2954 72
rect 2966 68 2970 72
rect 3038 68 3042 72
rect 2582 48 2586 52
rect 2598 48 2602 52
rect 2614 48 2618 52
rect 2838 48 2842 52
rect 2606 38 2610 42
rect 2862 38 2866 42
rect 2886 38 2890 42
rect 2566 18 2570 22
rect 2582 18 2586 22
rect 2678 18 2682 22
rect 2854 18 2858 22
rect 2538 3 2542 7
rect 2545 3 2549 7
rect 2702 8 2706 12
rect 2766 8 2770 12
rect 2862 8 2866 12
rect 2974 48 2978 52
rect 2950 38 2954 42
rect 2918 28 2922 32
rect 2966 28 2970 32
rect 3206 78 3210 82
rect 3310 318 3314 322
rect 3342 278 3346 282
rect 3358 318 3362 322
rect 3358 298 3362 302
rect 3318 258 3322 262
rect 3470 448 3474 452
rect 3510 388 3514 392
rect 3438 378 3442 382
rect 3486 368 3490 372
rect 3510 358 3514 362
rect 3462 348 3466 352
rect 3438 328 3442 332
rect 3390 308 3394 312
rect 3510 338 3514 342
rect 3446 298 3450 302
rect 3470 298 3474 302
rect 3414 268 3418 272
rect 3430 268 3434 272
rect 3278 248 3282 252
rect 3270 178 3274 182
rect 3246 158 3250 162
rect 3294 168 3298 172
rect 3398 238 3402 242
rect 3382 188 3386 192
rect 3390 168 3394 172
rect 3302 158 3306 162
rect 3318 158 3322 162
rect 3278 148 3282 152
rect 3286 148 3290 152
rect 3422 258 3426 262
rect 3454 258 3458 262
rect 3422 238 3426 242
rect 3414 218 3418 222
rect 3414 178 3418 182
rect 3430 168 3434 172
rect 3486 258 3490 262
rect 3478 248 3482 252
rect 3510 248 3514 252
rect 3470 198 3474 202
rect 3494 238 3498 242
rect 3542 568 3546 572
rect 3534 528 3538 532
rect 3542 508 3546 512
rect 3558 648 3562 652
rect 3534 468 3538 472
rect 3542 348 3546 352
rect 3542 288 3546 292
rect 3558 248 3562 252
rect 3542 208 3546 212
rect 3342 148 3346 152
rect 3382 148 3386 152
rect 3406 148 3410 152
rect 3550 158 3554 162
rect 3358 138 3362 142
rect 3382 138 3386 142
rect 3478 138 3482 142
rect 3286 128 3290 132
rect 3294 128 3298 132
rect 3326 128 3330 132
rect 3342 128 3346 132
rect 3366 128 3370 132
rect 3422 128 3426 132
rect 3454 128 3458 132
rect 3286 78 3290 82
rect 3134 68 3138 72
rect 3150 68 3154 72
rect 3206 68 3210 72
rect 3046 48 3050 52
rect 3134 48 3138 52
rect 3078 38 3082 42
rect 2982 18 2986 22
rect 3006 18 3010 22
rect 2910 8 2914 12
rect 3334 108 3338 112
rect 3310 98 3314 102
rect 3318 98 3322 102
rect 3374 108 3378 112
rect 3342 78 3346 82
rect 3486 118 3490 122
rect 3518 128 3522 132
rect 3430 98 3434 102
rect 3462 98 3466 102
rect 3510 98 3514 102
rect 3462 88 3466 92
rect 3478 78 3482 82
rect 3318 68 3322 72
rect 3334 68 3338 72
rect 3374 58 3378 62
rect 3534 58 3538 62
rect 3230 48 3234 52
rect 3158 38 3162 42
rect 3214 38 3218 42
rect 3310 28 3314 32
rect 3350 8 3354 12
<< metal3 >>
rect 992 3303 994 3307
rect 998 3303 1001 3307
rect 1006 3303 1008 3307
rect 2024 3303 2026 3307
rect 2030 3303 2033 3307
rect 2038 3303 2040 3307
rect 3040 3303 3042 3307
rect 3046 3303 3049 3307
rect 3054 3303 3056 3307
rect 690 3298 694 3301
rect 706 3298 734 3301
rect 1138 3298 1142 3301
rect 1290 3298 1294 3301
rect 1354 3298 1374 3301
rect 1410 3298 1414 3301
rect 1546 3298 1550 3301
rect 1650 3298 1654 3301
rect 1674 3298 1718 3301
rect 1730 3298 1734 3301
rect 1922 3298 1950 3301
rect 1994 3298 1998 3301
rect 2202 3298 2230 3301
rect 2258 3298 2262 3301
rect 2282 3298 2294 3301
rect 2466 3298 2470 3301
rect 2522 3298 2526 3301
rect 2634 3298 2638 3301
rect 2650 3298 2662 3301
rect 2810 3298 2814 3301
rect 2938 3298 2958 3301
rect 3082 3298 3086 3301
rect 606 3292 609 3298
rect 670 3292 673 3298
rect 1022 3292 1025 3298
rect 1054 3292 1057 3298
rect 1230 3292 1233 3298
rect 1598 3292 1601 3298
rect 2246 3292 2249 3298
rect 2926 3292 2929 3298
rect 786 3288 894 3291
rect 926 3288 934 3291
rect 938 3288 1014 3291
rect 1274 3288 1358 3291
rect 1642 3288 1670 3291
rect 1674 3288 2113 3291
rect 2122 3288 2158 3291
rect 2178 3288 2182 3291
rect 2234 3288 2238 3291
rect 2258 3288 2398 3291
rect 2470 3288 2478 3291
rect 2482 3288 2486 3291
rect 2630 3288 2646 3291
rect 2794 3288 2798 3291
rect 630 3282 633 3288
rect 114 3278 254 3281
rect 774 3281 777 3288
rect 730 3278 777 3281
rect 882 3278 886 3281
rect 906 3278 966 3281
rect 970 3278 1014 3281
rect 1026 3278 1086 3281
rect 1174 3278 1182 3281
rect 1186 3278 1534 3281
rect 1594 3278 1657 3281
rect 1654 3272 1657 3278
rect 1922 3278 2014 3281
rect 2018 3278 2070 3281
rect 2074 3278 2086 3281
rect 2110 3281 2113 3288
rect 2630 3282 2633 3288
rect 2110 3278 2142 3281
rect 2146 3278 2262 3281
rect 2402 3278 2502 3281
rect 2674 3278 2814 3281
rect 2818 3278 2950 3281
rect 2954 3278 2982 3281
rect 3122 3278 3126 3281
rect 3514 3278 3518 3281
rect 1702 3272 1705 3278
rect 322 3268 454 3271
rect 458 3268 478 3271
rect 690 3268 710 3271
rect 714 3268 718 3271
rect 746 3268 774 3271
rect 866 3268 1454 3271
rect 1490 3268 1518 3271
rect 1558 3268 1574 3271
rect 1642 3268 1646 3271
rect 1794 3268 2374 3271
rect 2378 3268 2454 3271
rect 2530 3268 2574 3271
rect 2638 3271 2641 3278
rect 3390 3272 3393 3278
rect 2638 3268 2694 3271
rect 3114 3268 3294 3271
rect 3314 3268 3318 3271
rect 3442 3268 3478 3271
rect 3514 3268 3518 3271
rect 94 3261 97 3268
rect 142 3261 145 3268
rect 94 3258 145 3261
rect 198 3261 201 3268
rect 198 3258 222 3261
rect 274 3258 334 3261
rect 354 3258 366 3261
rect 606 3261 609 3268
rect 606 3258 670 3261
rect 734 3261 737 3268
rect 1454 3262 1457 3268
rect 698 3258 737 3261
rect 770 3258 862 3261
rect 890 3258 910 3261
rect 930 3258 958 3261
rect 1010 3258 1038 3261
rect 1058 3258 1078 3261
rect 1106 3258 1190 3261
rect 1290 3258 1326 3261
rect 1362 3258 1374 3261
rect 1482 3258 1502 3261
rect 1558 3261 1561 3268
rect 1538 3258 1561 3261
rect 1570 3258 1702 3261
rect 1738 3258 1822 3261
rect 1842 3258 1846 3261
rect 1898 3259 1958 3261
rect 1898 3258 1961 3259
rect 2034 3258 2038 3261
rect 2042 3258 2054 3261
rect 2082 3258 2110 3261
rect 2146 3258 2158 3261
rect 2210 3258 2214 3261
rect 2306 3258 2310 3261
rect 2434 3258 2470 3261
rect 2514 3258 2558 3261
rect 2666 3258 2678 3261
rect 2706 3258 2758 3261
rect 2774 3261 2777 3268
rect 2854 3262 2857 3268
rect 3374 3262 3377 3268
rect 2774 3258 2798 3261
rect 2826 3258 2838 3261
rect 2922 3258 2942 3261
rect 3122 3258 3126 3261
rect 3178 3258 3182 3261
rect 3394 3258 3398 3261
rect 3402 3258 3438 3261
rect 3458 3258 3462 3261
rect 3510 3258 3518 3261
rect -26 3251 -22 3252
rect -26 3248 6 3251
rect 34 3248 158 3251
rect 162 3248 206 3251
rect 214 3248 342 3251
rect 358 3248 422 3251
rect 430 3251 433 3258
rect 430 3248 614 3251
rect 626 3248 790 3251
rect 886 3251 889 3258
rect 886 3248 942 3251
rect 1038 3251 1041 3258
rect 1246 3252 1249 3258
rect 1038 3248 1070 3251
rect 1082 3248 1118 3251
rect 1330 3248 1366 3251
rect 1370 3248 1422 3251
rect 1474 3248 1486 3251
rect 1510 3248 1638 3251
rect 1690 3248 1806 3251
rect 1810 3248 1878 3251
rect 1882 3248 1902 3251
rect 2230 3251 2233 3258
rect 3094 3252 3097 3258
rect 3366 3252 3369 3258
rect 2230 3248 2502 3251
rect 2530 3248 2590 3251
rect 2594 3248 2638 3251
rect 2846 3248 2854 3251
rect 2858 3248 2886 3251
rect 3010 3248 3054 3251
rect 3058 3248 3086 3251
rect 3370 3248 3398 3251
rect 3450 3248 3454 3251
rect 3498 3248 3550 3251
rect 214 3242 217 3248
rect 358 3242 361 3248
rect 474 3238 518 3241
rect 522 3238 550 3241
rect 554 3238 638 3241
rect 746 3238 870 3241
rect 874 3238 934 3241
rect 1022 3241 1025 3248
rect 1510 3242 1513 3248
rect 1022 3238 1054 3241
rect 1070 3238 1286 3241
rect 1298 3238 1401 3241
rect 1070 3232 1073 3238
rect 1398 3232 1401 3238
rect 1522 3238 1542 3241
rect 1578 3238 2198 3241
rect 2202 3238 2286 3241
rect 2442 3238 2614 3241
rect 2618 3238 2654 3241
rect 2730 3238 2830 3241
rect 2834 3238 3030 3241
rect 3034 3238 3070 3241
rect 3082 3238 3118 3241
rect 3146 3238 3294 3241
rect 3362 3238 3374 3241
rect 1430 3232 1433 3238
rect 178 3228 326 3231
rect 738 3228 750 3231
rect 1098 3228 1198 3231
rect 1770 3228 1934 3231
rect 2226 3228 2254 3231
rect 2786 3228 2894 3231
rect 3398 3231 3401 3238
rect 3398 3228 3470 3231
rect 3474 3228 3502 3231
rect 106 3218 126 3221
rect 138 3218 174 3221
rect 466 3218 654 3221
rect 658 3218 1078 3221
rect 1386 3218 1598 3221
rect 1858 3218 1950 3221
rect 2138 3218 2334 3221
rect 2338 3218 2358 3221
rect 2594 3218 2822 3221
rect 682 3208 910 3211
rect 1434 3208 1478 3211
rect 1882 3208 2446 3211
rect 2450 3208 2454 3211
rect 480 3203 482 3207
rect 486 3203 489 3207
rect 494 3203 496 3207
rect 1512 3203 1514 3207
rect 1518 3203 1521 3207
rect 1526 3203 1528 3207
rect 2536 3203 2538 3207
rect 2542 3203 2545 3207
rect 2550 3203 2552 3207
rect 1082 3198 1110 3201
rect 1266 3198 1502 3201
rect 1674 3198 1678 3201
rect 1962 3198 1974 3201
rect 3362 3198 3478 3201
rect 402 3188 494 3191
rect 1018 3188 1462 3191
rect 1466 3188 1678 3191
rect 3218 3188 3430 3191
rect 842 3178 998 3181
rect 1002 3178 1270 3181
rect 1402 3178 1510 3181
rect 1514 3178 1566 3181
rect 1874 3178 1958 3181
rect 1962 3178 2158 3181
rect 2970 3178 3102 3181
rect 3114 3178 3198 3181
rect 82 3168 86 3171
rect 322 3168 342 3171
rect 710 3171 713 3178
rect 1742 3172 1745 3178
rect 710 3168 734 3171
rect 738 3168 758 3171
rect 802 3168 822 3171
rect 834 3168 838 3171
rect 970 3168 1190 3171
rect 1206 3168 1246 3171
rect 1346 3168 1398 3171
rect 1602 3168 1686 3171
rect 1778 3168 1822 3171
rect 1858 3168 1902 3171
rect 1906 3168 2166 3171
rect 2170 3168 2230 3171
rect 2250 3168 2478 3171
rect 2482 3168 2486 3171
rect 2670 3171 2673 3178
rect 2670 3168 2702 3171
rect 2930 3168 3222 3171
rect 3226 3168 3230 3171
rect 3354 3168 3385 3171
rect 42 3158 46 3161
rect 122 3158 334 3161
rect 582 3161 585 3168
rect 578 3158 585 3161
rect 638 3161 641 3168
rect 1206 3162 1209 3168
rect 2710 3162 2713 3168
rect 3382 3162 3385 3168
rect 610 3158 641 3161
rect 722 3158 742 3161
rect 746 3158 785 3161
rect 794 3158 1022 3161
rect 1026 3158 1198 3161
rect 1310 3158 1382 3161
rect 1690 3158 1726 3161
rect 1938 3158 2030 3161
rect 2114 3158 2134 3161
rect 2226 3158 2294 3161
rect 2298 3158 2326 3161
rect 2338 3158 2422 3161
rect 2474 3158 2486 3161
rect 2506 3158 2646 3161
rect 2650 3158 2678 3161
rect 2962 3158 2974 3161
rect 3018 3158 3142 3161
rect 3218 3158 3270 3161
rect 3298 3158 3302 3161
rect 3338 3158 3358 3161
rect 3386 3158 3502 3161
rect 34 3148 94 3151
rect 138 3148 182 3151
rect 314 3148 318 3151
rect 506 3148 542 3151
rect 546 3148 598 3151
rect 642 3148 670 3151
rect 674 3148 774 3151
rect 782 3151 785 3158
rect 1286 3152 1289 3158
rect 1310 3152 1313 3158
rect 782 3148 806 3151
rect 810 3148 830 3151
rect 858 3148 862 3151
rect 906 3148 950 3151
rect 962 3148 1054 3151
rect 1066 3148 1110 3151
rect 1114 3148 1142 3151
rect 1146 3148 1158 3151
rect 1190 3148 1238 3151
rect 1258 3148 1281 3151
rect 1354 3148 1358 3151
rect 1374 3148 1462 3151
rect 1498 3148 1521 3151
rect 1674 3148 1694 3151
rect 1730 3148 1734 3151
rect 1770 3148 1782 3151
rect 1846 3151 1849 3158
rect 1826 3148 1849 3151
rect 1902 3151 1905 3158
rect 1866 3148 1905 3151
rect 1914 3148 1966 3151
rect 2018 3148 2054 3151
rect 18 3138 38 3141
rect 90 3138 134 3141
rect 154 3138 198 3141
rect 294 3141 297 3148
rect 1190 3142 1193 3148
rect 1278 3142 1281 3148
rect 1342 3142 1345 3148
rect 1374 3142 1377 3148
rect 1518 3142 1521 3148
rect 2066 3148 2150 3151
rect 2154 3148 2782 3151
rect 2890 3148 3246 3151
rect 3330 3148 3518 3151
rect 3590 3151 3594 3152
rect 3562 3148 3594 3151
rect 3038 3142 3041 3148
rect 3174 3142 3177 3148
rect 294 3138 414 3141
rect 530 3138 566 3141
rect 586 3138 606 3141
rect 666 3138 702 3141
rect 706 3138 766 3141
rect 786 3138 790 3141
rect 802 3138 974 3141
rect 994 3138 1062 3141
rect 1130 3138 1134 3141
rect 1138 3138 1166 3141
rect 1382 3138 1446 3141
rect 1650 3138 1670 3141
rect 1694 3138 1718 3141
rect 1738 3138 1974 3141
rect 2122 3138 2158 3141
rect 2306 3138 2310 3141
rect 2346 3138 2529 3141
rect 2538 3138 2574 3141
rect 2682 3138 2734 3141
rect 2778 3138 2782 3141
rect 3002 3138 3006 3141
rect 3326 3138 3358 3141
rect 3418 3138 3470 3141
rect 3498 3138 3534 3141
rect 26 3128 57 3131
rect 54 3122 57 3128
rect 118 3128 158 3131
rect 174 3128 206 3131
rect 282 3128 294 3131
rect 330 3128 366 3131
rect 370 3128 382 3131
rect 386 3128 462 3131
rect 610 3128 702 3131
rect 762 3128 806 3131
rect 810 3128 846 3131
rect 866 3128 966 3131
rect 970 3128 1070 3131
rect 1074 3128 1214 3131
rect 1382 3131 1385 3138
rect 1446 3132 1449 3138
rect 1694 3132 1697 3138
rect 2190 3132 2193 3138
rect 1242 3128 1385 3131
rect 1810 3128 1846 3131
rect 1850 3128 1870 3131
rect 2010 3128 2126 3131
rect 2170 3128 2174 3131
rect 2210 3128 2254 3131
rect 2258 3128 2262 3131
rect 2526 3131 2529 3138
rect 3326 3132 3329 3138
rect 2526 3128 2654 3131
rect 2658 3128 2686 3131
rect 2702 3128 2790 3131
rect 2802 3128 2806 3131
rect 3026 3128 3078 3131
rect 3386 3128 3398 3131
rect 118 3122 121 3128
rect 174 3122 177 3128
rect 146 3118 166 3121
rect 226 3118 310 3121
rect 450 3118 558 3121
rect 578 3118 686 3121
rect 690 3118 718 3121
rect 726 3121 729 3128
rect 1398 3122 1401 3128
rect 1662 3122 1665 3128
rect 726 3118 918 3121
rect 946 3118 974 3121
rect 978 3118 1014 3121
rect 1034 3118 1038 3121
rect 1098 3118 1102 3121
rect 1114 3118 1118 3121
rect 1138 3118 1182 3121
rect 1682 3118 1758 3121
rect 1882 3118 1990 3121
rect 2002 3118 2222 3121
rect 2454 3121 2457 3128
rect 2230 3118 2457 3121
rect 2470 3122 2473 3128
rect 2702 3122 2705 3128
rect 2514 3118 2526 3121
rect 2842 3118 2862 3121
rect 2874 3118 2918 3121
rect 2994 3118 3030 3121
rect 3034 3118 3094 3121
rect 3098 3118 3350 3121
rect 3386 3118 3462 3121
rect 602 3108 646 3111
rect 714 3108 750 3111
rect 754 3108 798 3111
rect 914 3108 918 3111
rect 1118 3111 1121 3118
rect 1118 3108 1294 3111
rect 1370 3108 1374 3111
rect 1650 3108 1806 3111
rect 1818 3108 1838 3111
rect 1842 3108 1966 3111
rect 2138 3108 2206 3111
rect 2230 3111 2233 3118
rect 2218 3108 2233 3111
rect 2370 3108 2374 3111
rect 2394 3108 2582 3111
rect 2690 3108 2750 3111
rect 3178 3108 3182 3111
rect 3186 3108 3238 3111
rect 3306 3108 3422 3111
rect 992 3103 994 3107
rect 998 3103 1001 3107
rect 1006 3103 1008 3107
rect 2024 3103 2026 3107
rect 2030 3103 2033 3107
rect 2038 3103 2040 3107
rect 3040 3103 3042 3107
rect 3046 3103 3049 3107
rect 3054 3103 3056 3107
rect 570 3098 774 3101
rect 778 3098 814 3101
rect 850 3098 862 3101
rect 922 3098 966 3101
rect 1018 3098 1230 3101
rect 1258 3098 1462 3101
rect 1546 3098 1654 3101
rect 1658 3098 1766 3101
rect 1834 3098 1894 3101
rect 2050 3098 2166 3101
rect 2170 3098 2270 3101
rect 2466 3098 2510 3101
rect 58 3088 78 3091
rect 290 3088 358 3091
rect 606 3088 614 3091
rect 822 3088 830 3091
rect 834 3088 870 3091
rect 1134 3088 1158 3091
rect 1330 3088 1406 3091
rect 1434 3088 1526 3091
rect 1574 3088 1582 3091
rect 1586 3088 1622 3091
rect 1642 3088 1662 3091
rect 1814 3088 1862 3091
rect 1954 3088 1990 3091
rect 2010 3088 2014 3091
rect 2146 3088 2214 3091
rect 2250 3088 2286 3091
rect 2322 3088 2494 3091
rect 3090 3088 3174 3091
rect 3322 3088 3334 3091
rect 42 3078 62 3081
rect 66 3078 134 3081
rect 322 3078 350 3081
rect 598 3081 601 3088
rect 474 3078 601 3081
rect 610 3078 622 3081
rect 682 3078 846 3081
rect 850 3078 902 3081
rect 958 3081 961 3088
rect 1134 3082 1137 3088
rect 922 3078 961 3081
rect 1082 3078 1102 3081
rect 1130 3078 1134 3081
rect 1146 3078 1150 3081
rect 1210 3078 1214 3081
rect 1290 3078 1294 3081
rect 1298 3078 1374 3081
rect 1514 3078 1590 3081
rect 1710 3081 1713 3088
rect 1626 3078 1713 3081
rect 1814 3082 1817 3088
rect 1930 3078 2065 3081
rect 2062 3072 2065 3078
rect 2162 3078 2166 3081
rect 2186 3078 2222 3081
rect 2230 3081 2233 3088
rect 2230 3078 2262 3081
rect 2434 3078 2438 3081
rect 2450 3078 2470 3081
rect 2522 3078 2534 3081
rect 2858 3078 2862 3081
rect 2866 3078 2990 3081
rect 3214 3081 3217 3088
rect 3214 3078 3342 3081
rect 2086 3072 2089 3078
rect 2094 3072 2097 3078
rect 10 3068 38 3071
rect 70 3068 78 3071
rect 82 3068 166 3071
rect 178 3068 190 3071
rect 210 3068 238 3071
rect 242 3068 398 3071
rect 402 3068 478 3071
rect 482 3068 582 3071
rect 586 3068 1614 3071
rect 1626 3068 1630 3071
rect 1682 3068 1750 3071
rect 1826 3068 1830 3071
rect 1834 3068 1886 3071
rect 1922 3068 2006 3071
rect 2114 3068 2150 3071
rect 2178 3068 2182 3071
rect 2390 3071 2393 3078
rect 2290 3068 2393 3071
rect 2410 3068 2462 3071
rect 2466 3068 2486 3071
rect 2514 3068 2558 3071
rect 2586 3068 2654 3071
rect 2702 3071 2705 3078
rect 2658 3068 2705 3071
rect 2786 3068 3166 3071
rect 3170 3068 3254 3071
rect 34 3058 142 3061
rect 202 3058 206 3061
rect 210 3058 246 3061
rect 338 3058 342 3061
rect 450 3058 462 3061
rect 562 3059 566 3061
rect 558 3058 566 3059
rect 602 3058 614 3061
rect 762 3058 806 3061
rect 810 3058 854 3061
rect 858 3058 918 3061
rect 970 3058 1022 3061
rect 1054 3058 1062 3061
rect 1066 3058 1118 3061
rect 1122 3058 1142 3061
rect 1338 3058 1702 3061
rect 1706 3058 1782 3061
rect 1790 3061 1793 3068
rect 1790 3058 2062 3061
rect 2074 3058 2102 3061
rect 2186 3058 2206 3061
rect 2346 3058 2350 3061
rect 2426 3058 2494 3061
rect 2514 3058 2521 3061
rect 2626 3058 2721 3061
rect 2786 3058 2806 3061
rect 2822 3058 2846 3061
rect 2914 3058 2918 3061
rect 2954 3058 2990 3061
rect 3050 3058 3062 3061
rect 3074 3059 3126 3061
rect 3074 3058 3129 3059
rect 3218 3058 3249 3061
rect 2126 3052 2129 3058
rect -26 3051 -22 3052
rect -26 3048 6 3051
rect 10 3048 78 3051
rect 202 3048 222 3051
rect 226 3048 254 3051
rect 258 3048 286 3051
rect 338 3048 342 3051
rect 434 3048 470 3051
rect 546 3048 590 3051
rect 594 3048 622 3051
rect 798 3048 942 3051
rect 1042 3048 1089 3051
rect 1130 3048 1246 3051
rect 1274 3048 1310 3051
rect 1370 3048 1398 3051
rect 1418 3048 1446 3051
rect 1474 3048 1478 3051
rect 1490 3048 1494 3051
rect 1554 3048 1582 3051
rect 1586 3048 1630 3051
rect 1658 3048 1902 3051
rect 1906 3048 1982 3051
rect 1994 3048 2014 3051
rect 2106 3048 2118 3051
rect 2422 3051 2425 3058
rect 2518 3052 2521 3058
rect 2718 3052 2721 3058
rect 2822 3052 2825 3058
rect 3246 3052 3249 3058
rect 2202 3048 2417 3051
rect 2422 3048 2454 3051
rect 2490 3048 2502 3051
rect 2594 3048 2630 3051
rect 3074 3048 3086 3051
rect 3130 3048 3190 3051
rect 798 3042 801 3048
rect 90 3038 118 3041
rect 122 3038 209 3041
rect 206 3032 209 3038
rect 238 3038 270 3041
rect 362 3038 382 3041
rect 602 3038 606 3041
rect 950 3041 953 3048
rect 1086 3042 1089 3048
rect 950 3038 1078 3041
rect 1122 3038 1134 3041
rect 1226 3038 1313 3041
rect 1322 3038 1430 3041
rect 1434 3038 1566 3041
rect 1614 3038 1622 3041
rect 1626 3038 1646 3041
rect 1694 3038 1734 3041
rect 1850 3038 1862 3041
rect 1866 3038 1950 3041
rect 1978 3038 2046 3041
rect 2050 3038 2190 3041
rect 2194 3038 2262 3041
rect 2266 3038 2302 3041
rect 2306 3038 2318 3041
rect 2414 3041 2417 3048
rect 2414 3038 2430 3041
rect 2450 3038 2510 3041
rect 2514 3038 2670 3041
rect 2674 3038 2718 3041
rect 2770 3038 3006 3041
rect 3202 3038 3222 3041
rect 3322 3038 3334 3041
rect 238 3032 241 3038
rect 1310 3032 1313 3038
rect 458 3028 542 3031
rect 594 3028 686 3031
rect 690 3028 694 3031
rect 698 3028 726 3031
rect 834 3028 1118 3031
rect 1378 3028 1438 3031
rect 1694 3031 1697 3038
rect 1442 3028 1697 3031
rect 1862 3028 1902 3031
rect 1906 3028 1982 3031
rect 2082 3028 2110 3031
rect 2114 3028 2158 3031
rect 2162 3028 2206 3031
rect 2450 3028 2518 3031
rect 2530 3028 3054 3031
rect 1702 3022 1705 3028
rect 1862 3022 1865 3028
rect 522 3018 718 3021
rect 738 3018 934 3021
rect 938 3018 1038 3021
rect 1042 3018 1046 3021
rect 1098 3018 1222 3021
rect 1314 3018 1390 3021
rect 1426 3018 1478 3021
rect 1554 3018 1582 3021
rect 2274 3018 2574 3021
rect 2762 3018 2830 3021
rect 1230 3012 1233 3018
rect 714 3008 734 3011
rect 914 3008 1150 3011
rect 1306 3008 1502 3011
rect 1730 3008 2438 3011
rect 2562 3008 2806 3011
rect 2810 3008 3310 3011
rect 480 3003 482 3007
rect 486 3003 489 3007
rect 494 3003 496 3007
rect 1512 3003 1514 3007
rect 1518 3003 1521 3007
rect 1526 3003 1528 3007
rect 2536 3003 2538 3007
rect 2542 3003 2545 3007
rect 2550 3003 2552 3007
rect 674 2998 734 3001
rect 762 2998 830 3001
rect 1090 2998 1102 3001
rect 1346 2998 1430 3001
rect 1474 2998 1478 3001
rect 1498 2998 1502 3001
rect 1570 2998 1822 3001
rect 1834 2998 2214 3001
rect 2434 2998 2470 3001
rect 2714 2998 2782 3001
rect 2986 2998 2990 3001
rect 730 2988 854 2991
rect 938 2988 974 2991
rect 1058 2988 1238 2991
rect 1250 2988 1254 2991
rect 1430 2991 1433 2998
rect 2238 2992 2241 2998
rect 1430 2988 1558 2991
rect 1594 2988 1774 2991
rect 1842 2988 1886 2991
rect 2982 2988 3006 2991
rect 2982 2982 2985 2988
rect 418 2978 654 2981
rect 722 2978 886 2981
rect 890 2978 918 2981
rect 922 2978 926 2981
rect 930 2978 942 2981
rect 1226 2978 1353 2981
rect 1362 2978 1454 2981
rect 1466 2978 1774 2981
rect 1842 2978 1870 2981
rect 2050 2978 2230 2981
rect 2242 2978 2246 2981
rect 2442 2978 2734 2981
rect 3026 2978 3078 2981
rect 3514 2978 3518 2981
rect 1350 2972 1353 2978
rect 106 2968 110 2971
rect 858 2968 1118 2971
rect 1186 2968 1230 2971
rect 1370 2968 1470 2971
rect 1482 2968 1726 2971
rect 1730 2968 1742 2971
rect 1862 2968 1894 2971
rect 1990 2971 1993 2978
rect 1990 2968 2062 2971
rect 3490 2968 3518 2971
rect 26 2958 86 2961
rect 138 2958 182 2961
rect 186 2958 190 2961
rect 194 2958 254 2961
rect 282 2958 286 2961
rect 378 2958 390 2961
rect 670 2961 673 2968
rect 670 2958 710 2961
rect 730 2958 782 2961
rect 850 2958 870 2961
rect 954 2958 1022 2961
rect 1098 2958 1118 2961
rect 1146 2958 1158 2961
rect 1162 2958 1214 2961
rect 1318 2961 1321 2968
rect 1862 2962 1865 2968
rect 1218 2958 1321 2961
rect 1362 2958 1414 2961
rect 1418 2958 1430 2961
rect 1442 2958 1446 2961
rect 1458 2958 1494 2961
rect 1506 2958 1518 2961
rect 1538 2958 1686 2961
rect 1738 2958 1782 2961
rect 1890 2958 2046 2961
rect 2074 2958 2150 2961
rect 2174 2961 2177 2968
rect 2174 2958 2182 2961
rect 2210 2958 2278 2961
rect 2462 2961 2465 2968
rect 2338 2958 2465 2961
rect 2522 2958 2558 2961
rect 2934 2961 2937 2968
rect 2966 2961 2969 2968
rect 3542 2962 3545 2968
rect 2842 2958 2873 2961
rect 2934 2958 2969 2961
rect 2986 2958 3014 2961
rect 3018 2958 3206 2961
rect 3250 2958 3262 2961
rect 3274 2958 3278 2961
rect 1062 2952 1065 2958
rect 2870 2952 2873 2958
rect 42 2948 62 2951
rect 66 2948 150 2951
rect 234 2948 238 2951
rect 266 2948 270 2951
rect 346 2948 366 2951
rect 434 2948 534 2951
rect 626 2948 630 2951
rect 634 2948 670 2951
rect 698 2948 734 2951
rect 746 2948 822 2951
rect 850 2948 854 2951
rect 858 2948 1014 2951
rect 1098 2948 1694 2951
rect 1698 2948 2046 2951
rect 2066 2948 2086 2951
rect 2114 2948 2134 2951
rect 2178 2948 2182 2951
rect 2202 2948 2222 2951
rect 2274 2948 2326 2951
rect 2498 2948 2526 2951
rect 2530 2948 2542 2951
rect 2546 2948 2582 2951
rect 2586 2948 2662 2951
rect 2882 2948 2894 2951
rect 2922 2948 2942 2951
rect 3018 2948 3046 2951
rect 3090 2948 3102 2951
rect 3106 2948 3110 2951
rect 3162 2948 3193 2951
rect 3234 2948 3254 2951
rect 3258 2948 3302 2951
rect 3474 2948 3486 2951
rect 3490 2948 3534 2951
rect 3538 2948 3542 2951
rect 1014 2942 1017 2948
rect 1046 2942 1049 2948
rect 2366 2942 2369 2948
rect 3190 2942 3193 2948
rect 50 2938 86 2941
rect 90 2938 126 2941
rect 210 2938 230 2941
rect 314 2938 334 2941
rect 354 2938 390 2941
rect 394 2938 406 2941
rect 474 2938 558 2941
rect 618 2938 678 2941
rect 682 2938 742 2941
rect 810 2938 814 2941
rect 994 2938 998 2941
rect 1082 2938 1102 2941
rect 1130 2938 1134 2941
rect 1194 2938 1222 2941
rect 1234 2938 1254 2941
rect 1282 2938 1310 2941
rect 1314 2938 1326 2941
rect 1330 2938 1574 2941
rect 1578 2938 1633 2941
rect 42 2928 54 2931
rect 82 2928 102 2931
rect 178 2928 198 2931
rect 346 2928 430 2931
rect 434 2928 438 2931
rect 578 2928 582 2931
rect 618 2928 630 2931
rect 690 2928 766 2931
rect 790 2931 793 2938
rect 778 2928 793 2931
rect 802 2928 806 2931
rect 834 2928 841 2931
rect 898 2928 910 2931
rect 926 2931 929 2938
rect 922 2928 929 2931
rect 966 2932 969 2938
rect 974 2932 977 2938
rect 1010 2928 1046 2931
rect 1050 2928 1070 2931
rect 1174 2931 1177 2938
rect 1630 2932 1633 2938
rect 1826 2938 1830 2941
rect 1858 2938 1878 2941
rect 1898 2938 1918 2941
rect 1994 2938 1998 2941
rect 2034 2938 2078 2941
rect 2082 2938 2214 2941
rect 2226 2938 2270 2941
rect 2282 2938 2310 2941
rect 2506 2938 2510 2941
rect 2738 2938 2878 2941
rect 2914 2938 2934 2941
rect 3042 2938 3062 2941
rect 3066 2938 3078 2941
rect 3138 2938 3150 2941
rect 1766 2932 1769 2938
rect 1878 2932 1881 2938
rect 1934 2932 1937 2938
rect 2014 2932 2017 2938
rect 1106 2928 1177 2931
rect 1186 2928 1214 2931
rect 1226 2928 1262 2931
rect 1326 2928 1342 2931
rect 1354 2928 1358 2931
rect 1442 2928 1454 2931
rect 1510 2928 1598 2931
rect 1650 2928 1654 2931
rect 1794 2928 1798 2931
rect 1866 2928 1870 2931
rect 2018 2928 2070 2931
rect 2082 2928 2438 2931
rect 2466 2928 2494 2931
rect 2506 2928 2606 2931
rect 2674 2928 2694 2931
rect 2698 2928 2798 2931
rect 2938 2928 2942 2931
rect 3102 2931 3105 2938
rect 3102 2928 3142 2931
rect 3178 2928 3206 2931
rect 3210 2928 3254 2931
rect 3274 2928 3278 2931
rect 3294 2931 3297 2938
rect 3374 2931 3377 2938
rect 3282 2928 3377 2931
rect 3422 2932 3425 2938
rect 14 2918 22 2921
rect 26 2918 46 2921
rect 58 2918 134 2921
rect 138 2918 198 2921
rect 234 2918 414 2921
rect 698 2918 718 2921
rect 862 2921 865 2928
rect 1326 2922 1329 2928
rect 1510 2922 1513 2928
rect 1622 2922 1625 2928
rect 762 2918 865 2921
rect 870 2918 1046 2921
rect 1254 2918 1318 2921
rect 1354 2918 1374 2921
rect 1378 2918 1382 2921
rect 1426 2918 1510 2921
rect 1554 2918 1606 2921
rect 1658 2918 1734 2921
rect 1742 2921 1745 2928
rect 1742 2918 1806 2921
rect 1898 2918 1990 2921
rect 2014 2918 2094 2921
rect 2098 2918 2126 2921
rect 2378 2918 2478 2921
rect 2718 2918 2726 2921
rect 2730 2918 2862 2921
rect 3058 2918 3113 2921
rect 3122 2918 3126 2921
rect 3162 2918 3198 2921
rect 3274 2918 3350 2921
rect 138 2908 142 2911
rect 154 2908 238 2911
rect 298 2908 446 2911
rect 450 2908 478 2911
rect 482 2908 646 2911
rect 870 2911 873 2918
rect 650 2908 873 2911
rect 1026 2908 1038 2911
rect 1254 2911 1257 2918
rect 1162 2908 1257 2911
rect 1266 2908 1406 2911
rect 1418 2908 1566 2911
rect 1570 2908 1606 2911
rect 1618 2908 1646 2911
rect 1722 2908 1838 2911
rect 1874 2908 1910 2911
rect 2014 2911 2017 2918
rect 1922 2908 2017 2911
rect 2122 2908 2150 2911
rect 2154 2908 2446 2911
rect 2778 2908 2814 2911
rect 2818 2908 2854 2911
rect 3110 2911 3113 2918
rect 3110 2908 3182 2911
rect 3186 2908 3214 2911
rect 3218 2908 3246 2911
rect 3370 2908 3398 2911
rect 992 2903 994 2907
rect 998 2903 1001 2907
rect 1006 2903 1008 2907
rect 114 2898 214 2901
rect 218 2898 262 2901
rect 282 2898 302 2901
rect 410 2898 414 2901
rect 450 2898 454 2901
rect 658 2898 966 2901
rect 1034 2898 1086 2901
rect 1114 2898 1118 2901
rect 1154 2898 1438 2901
rect 1458 2898 1470 2901
rect 1614 2901 1617 2908
rect 2024 2903 2026 2907
rect 2030 2903 2033 2907
rect 2038 2903 2040 2907
rect 3040 2903 3042 2907
rect 3046 2903 3049 2907
rect 3054 2903 3056 2907
rect 3534 2902 3537 2908
rect 1474 2898 1617 2901
rect 1818 2898 1822 2901
rect 1842 2898 1926 2901
rect 1938 2898 1982 2901
rect 2106 2898 2230 2901
rect 2290 2898 2318 2901
rect 2474 2898 2502 2901
rect 2650 2898 2774 2901
rect 2778 2898 2822 2901
rect 3442 2898 3457 2901
rect 3522 2898 3526 2901
rect 74 2888 190 2891
rect 194 2888 286 2891
rect 346 2888 462 2891
rect 634 2888 726 2891
rect 730 2888 830 2891
rect 842 2888 854 2891
rect 954 2888 982 2891
rect 1074 2888 1078 2891
rect 1114 2888 1118 2891
rect 1138 2888 1142 2891
rect 1170 2888 1262 2891
rect 1306 2888 1566 2891
rect 1586 2888 2150 2891
rect 2154 2888 2238 2891
rect 2246 2888 2254 2891
rect 2258 2888 2302 2891
rect 2306 2888 2390 2891
rect 2402 2888 2462 2891
rect 2490 2888 2502 2891
rect 2506 2888 2534 2891
rect 2634 2888 2694 2891
rect 2754 2888 2926 2891
rect 3078 2888 3086 2891
rect 3090 2888 3118 2891
rect 3122 2888 3198 2891
rect 3378 2888 3446 2891
rect 3454 2891 3457 2898
rect 3454 2888 3537 2891
rect 10 2878 97 2881
rect 162 2878 238 2881
rect 250 2878 278 2881
rect 294 2881 297 2888
rect 294 2878 318 2881
rect 402 2878 422 2881
rect 470 2881 473 2888
rect 1054 2882 1057 2888
rect 458 2878 473 2881
rect 554 2878 558 2881
rect 578 2878 662 2881
rect 674 2878 686 2881
rect 738 2878 782 2881
rect 826 2878 878 2881
rect 882 2878 902 2881
rect 938 2878 1030 2881
rect 1066 2878 1206 2881
rect 1210 2878 1230 2881
rect 1242 2878 1262 2881
rect 1278 2881 1281 2888
rect 1266 2878 1281 2881
rect 1290 2878 1462 2881
rect 1466 2878 1478 2881
rect 1546 2878 1550 2881
rect 1558 2878 1630 2881
rect 1634 2878 1662 2881
rect 1730 2878 1750 2881
rect 1770 2878 1822 2881
rect 1850 2878 1854 2881
rect 1874 2878 1886 2881
rect 1970 2878 1982 2881
rect 1986 2878 2110 2881
rect 2122 2878 2206 2881
rect 2218 2878 2358 2881
rect 2398 2881 2401 2888
rect 2398 2878 2430 2881
rect 2458 2878 2590 2881
rect 2610 2878 2638 2881
rect 2730 2878 2758 2881
rect 2762 2878 2782 2881
rect 2786 2878 2886 2881
rect 3018 2878 3054 2881
rect 3058 2878 3078 2881
rect 3122 2878 3182 2881
rect 3210 2878 3230 2881
rect 3322 2878 3326 2881
rect 3338 2878 3342 2881
rect 3350 2881 3353 2888
rect 3534 2882 3537 2888
rect 3350 2878 3374 2881
rect 3438 2878 3478 2881
rect 3490 2878 3494 2881
rect 3514 2878 3518 2881
rect 94 2872 97 2878
rect -26 2871 -22 2872
rect -26 2868 22 2871
rect 26 2868 86 2871
rect 154 2868 174 2871
rect 242 2868 334 2871
rect 338 2868 350 2871
rect 370 2868 374 2871
rect 426 2868 430 2871
rect 466 2868 638 2871
rect 642 2868 654 2871
rect 730 2868 734 2871
rect 762 2868 766 2871
rect 862 2868 886 2871
rect 906 2868 910 2871
rect 938 2868 942 2871
rect 986 2868 1062 2871
rect 1074 2868 1094 2871
rect 1138 2868 1145 2871
rect 1186 2868 1286 2871
rect 1378 2868 1382 2871
rect 1386 2868 1398 2871
rect 1434 2868 1478 2871
rect 1558 2871 1561 2878
rect 3438 2872 3441 2878
rect 1482 2868 1561 2871
rect 1578 2868 1622 2871
rect 1658 2868 1718 2871
rect 1730 2868 1734 2871
rect 1778 2868 2150 2871
rect 2170 2868 2198 2871
rect 2250 2868 2254 2871
rect 2258 2868 2286 2871
rect 2334 2868 2374 2871
rect 2378 2868 2414 2871
rect 2426 2868 2446 2871
rect 2474 2868 2478 2871
rect 2490 2868 2494 2871
rect 2530 2868 2574 2871
rect 2602 2868 2670 2871
rect 2690 2868 2710 2871
rect 2994 2868 2998 2871
rect 3074 2868 3102 2871
rect 3106 2868 3126 2871
rect 3250 2868 3326 2871
rect 3330 2868 3350 2871
rect 3370 2868 3414 2871
rect 3482 2868 3502 2871
rect 3530 2868 3534 2871
rect 34 2858 38 2861
rect 86 2861 89 2868
rect 110 2861 113 2868
rect 86 2858 113 2861
rect 130 2858 206 2861
rect 250 2858 390 2861
rect 514 2858 518 2861
rect 602 2858 638 2861
rect 642 2858 718 2861
rect 774 2861 777 2868
rect 722 2858 777 2861
rect 814 2861 817 2868
rect 862 2862 865 2868
rect 1142 2862 1145 2868
rect 2334 2862 2337 2868
rect 2790 2862 2793 2868
rect 794 2858 817 2861
rect 850 2858 854 2861
rect 970 2858 1126 2861
rect 1178 2858 1302 2861
rect 1330 2858 1374 2861
rect 1378 2858 1382 2861
rect 1482 2858 1486 2861
rect 1506 2858 1638 2861
rect 1738 2858 1782 2861
rect 1842 2858 1846 2861
rect 1858 2858 1902 2861
rect 1922 2858 1926 2861
rect 1930 2858 1950 2861
rect 1994 2858 1998 2861
rect 2066 2858 2078 2861
rect 2218 2858 2222 2861
rect 2226 2858 2238 2861
rect 2274 2858 2286 2861
rect 2298 2858 2334 2861
rect 2362 2858 2494 2861
rect 2498 2858 2550 2861
rect 2570 2858 2598 2861
rect 2642 2858 2702 2861
rect 2730 2858 2766 2861
rect 2818 2858 2822 2861
rect 2826 2858 2878 2861
rect 3002 2858 3182 2861
rect 3186 2858 3198 2861
rect 3266 2858 3326 2861
rect 3330 2858 3342 2861
rect 3346 2858 3350 2861
rect 3474 2858 3494 2861
rect 3530 2858 3542 2861
rect -26 2851 -22 2852
rect -26 2848 6 2851
rect 18 2848 70 2851
rect 106 2848 110 2851
rect 210 2848 270 2851
rect 274 2848 294 2851
rect 314 2848 326 2851
rect 362 2848 366 2851
rect 410 2848 454 2851
rect 466 2848 486 2851
rect 602 2848 614 2851
rect 690 2848 710 2851
rect 1034 2848 1081 2851
rect 1146 2848 1174 2851
rect 1202 2848 1222 2851
rect 1226 2848 1230 2851
rect 1274 2848 1310 2851
rect 1330 2848 1382 2851
rect 1386 2848 1390 2851
rect 1410 2848 1526 2851
rect 1614 2848 1654 2851
rect 1662 2848 1694 2851
rect 1722 2848 1750 2851
rect 1770 2848 1774 2851
rect 1786 2848 1790 2851
rect 1818 2848 1902 2851
rect 1938 2848 1942 2851
rect 1954 2848 1958 2851
rect 1962 2848 1966 2851
rect 2058 2848 2118 2851
rect 2210 2848 2270 2851
rect 2330 2848 2366 2851
rect 2446 2848 2454 2851
rect 2458 2848 2470 2851
rect 2578 2848 2582 2851
rect 2690 2848 2742 2851
rect 2770 2848 2790 2851
rect 2802 2848 2806 2851
rect 3026 2848 3086 2851
rect 3090 2848 3113 2851
rect 3266 2848 3294 2851
rect 3314 2848 3334 2851
rect 3446 2851 3449 2858
rect 3446 2848 3510 2851
rect 50 2838 150 2841
rect 302 2841 305 2848
rect 1078 2842 1081 2848
rect 1614 2842 1617 2848
rect 1662 2842 1665 2848
rect 302 2838 582 2841
rect 586 2838 622 2841
rect 674 2838 910 2841
rect 1202 2838 1270 2841
rect 1290 2838 1374 2841
rect 1410 2838 1414 2841
rect 1434 2838 1590 2841
rect 1754 2838 1806 2841
rect 1966 2841 1969 2848
rect 1966 2838 2198 2841
rect 2410 2838 2494 2841
rect 2662 2841 2665 2848
rect 3110 2842 3113 2848
rect 3350 2842 3353 2848
rect 2662 2838 2670 2841
rect 2746 2838 2846 2841
rect 2930 2838 3094 2841
rect 3138 2838 3286 2841
rect 3318 2838 3334 2841
rect 98 2828 134 2831
rect 282 2828 286 2831
rect 410 2828 430 2831
rect 482 2828 526 2831
rect 622 2831 625 2838
rect 622 2828 718 2831
rect 926 2831 929 2838
rect 3318 2832 3321 2838
rect 730 2828 929 2831
rect 954 2828 1030 2831
rect 1074 2828 1702 2831
rect 1706 2828 1830 2831
rect 1906 2828 1982 2831
rect 1986 2828 2006 2831
rect 2010 2828 2094 2831
rect 2098 2828 2142 2831
rect 2162 2828 2182 2831
rect 2194 2828 2206 2831
rect 2442 2828 2614 2831
rect 2738 2828 2806 2831
rect 106 2818 118 2821
rect 430 2821 433 2828
rect 430 2818 782 2821
rect 850 2818 870 2821
rect 874 2818 1118 2821
rect 1250 2818 1702 2821
rect 1706 2818 1958 2821
rect 1970 2818 2137 2821
rect 2162 2818 2302 2821
rect 2326 2821 2329 2828
rect 2326 2818 2478 2821
rect 2490 2818 2694 2821
rect 2970 2818 2982 2821
rect 3174 2821 3177 2828
rect 3174 2818 3206 2821
rect 3322 2818 3326 2821
rect 34 2808 166 2811
rect 546 2808 654 2811
rect 666 2808 726 2811
rect 970 2808 1110 2811
rect 1138 2808 1318 2811
rect 1354 2808 1390 2811
rect 1594 2808 1598 2811
rect 1642 2808 1646 2811
rect 1674 2808 1678 2811
rect 1730 2808 1774 2811
rect 2026 2808 2126 2811
rect 2134 2811 2137 2818
rect 2134 2808 2486 2811
rect 3154 2808 3158 2811
rect 3162 2808 3174 2811
rect 3178 2808 3214 2811
rect 3290 2808 3446 2811
rect 480 2803 482 2807
rect 486 2803 489 2807
rect 494 2803 496 2807
rect 1512 2803 1514 2807
rect 1518 2803 1521 2807
rect 1526 2803 1528 2807
rect 1806 2802 1809 2808
rect 2536 2803 2538 2807
rect 2542 2803 2545 2807
rect 2550 2803 2552 2807
rect 2574 2802 2577 2808
rect 378 2798 470 2801
rect 562 2798 590 2801
rect 642 2798 678 2801
rect 690 2798 798 2801
rect 818 2798 1134 2801
rect 1138 2798 1150 2801
rect 1274 2798 1358 2801
rect 1930 2798 2174 2801
rect 2186 2798 2222 2801
rect 2250 2798 2366 2801
rect 2594 2798 2974 2801
rect 3034 2798 3406 2801
rect 806 2792 809 2798
rect 3454 2792 3457 2798
rect 386 2788 566 2791
rect 586 2788 622 2791
rect 626 2788 686 2791
rect 834 2788 990 2791
rect 1094 2788 1102 2791
rect 1106 2788 1110 2791
rect 1122 2788 1286 2791
rect 1294 2788 1302 2791
rect 1306 2788 1406 2791
rect 1530 2788 1542 2791
rect 1578 2788 2446 2791
rect 2498 2788 2569 2791
rect 3090 2788 3334 2791
rect 2566 2782 2569 2788
rect 3478 2782 3481 2788
rect 266 2778 390 2781
rect 394 2778 886 2781
rect 890 2778 910 2781
rect 914 2778 1046 2781
rect 1050 2778 1350 2781
rect 1498 2778 1726 2781
rect 1738 2778 1974 2781
rect 2042 2778 2246 2781
rect 2274 2778 2374 2781
rect 2378 2778 2422 2781
rect 2426 2778 2430 2781
rect 2690 2778 2710 2781
rect 2762 2778 2806 2781
rect 3010 2778 3254 2781
rect 3322 2778 3470 2781
rect 1574 2772 1577 2778
rect 138 2768 398 2771
rect 402 2768 622 2771
rect 642 2768 790 2771
rect 794 2768 822 2771
rect 826 2768 934 2771
rect 946 2768 950 2771
rect 962 2768 1238 2771
rect 1242 2768 1534 2771
rect 1546 2768 1550 2771
rect 1698 2768 1790 2771
rect 1810 2768 1822 2771
rect 1866 2768 1870 2771
rect 1874 2768 1926 2771
rect 2002 2768 2102 2771
rect 2110 2768 2118 2771
rect 2122 2768 2166 2771
rect 2194 2768 2254 2771
rect 2266 2768 2502 2771
rect 2602 2768 2926 2771
rect 3018 2768 3022 2771
rect 3114 2768 3182 2771
rect 3186 2768 3222 2771
rect 3226 2768 3262 2771
rect 3434 2768 3478 2771
rect 3490 2768 3502 2771
rect 3534 2771 3537 2778
rect 3506 2768 3537 2771
rect 90 2758 166 2761
rect 170 2758 174 2761
rect 270 2758 278 2761
rect 282 2758 302 2761
rect 434 2758 446 2761
rect 450 2758 846 2761
rect 858 2758 862 2761
rect 882 2758 942 2761
rect 1018 2758 1102 2761
rect 1114 2758 1150 2761
rect 1202 2758 1214 2761
rect 1258 2758 1374 2761
rect 1378 2758 1398 2761
rect 1458 2758 1462 2761
rect 1546 2758 1598 2761
rect 1694 2761 1697 2768
rect 1634 2758 1697 2761
rect 1706 2758 1742 2761
rect 1794 2758 1854 2761
rect 1858 2758 1878 2761
rect 1954 2758 2046 2761
rect 2058 2758 2062 2761
rect 2090 2758 2166 2761
rect 2182 2758 2257 2761
rect 2266 2758 2278 2761
rect 2450 2758 2462 2761
rect 2530 2758 2550 2761
rect 2554 2758 2558 2761
rect 2674 2758 2734 2761
rect 2738 2758 2798 2761
rect 2926 2761 2929 2768
rect 2890 2758 2929 2761
rect 3074 2758 3134 2761
rect 3170 2758 3174 2761
rect 3194 2758 3198 2761
rect 3242 2758 3278 2761
rect 3362 2758 3526 2761
rect 1230 2752 1233 2758
rect 2182 2752 2185 2758
rect 34 2748 54 2751
rect 154 2748 166 2751
rect 258 2748 286 2751
rect 290 2748 310 2751
rect 330 2748 334 2751
rect 378 2748 438 2751
rect 466 2748 486 2751
rect 514 2748 542 2751
rect 554 2748 558 2751
rect 586 2748 662 2751
rect 666 2748 702 2751
rect 766 2748 870 2751
rect 954 2748 990 2751
rect 1090 2748 1126 2751
rect 1178 2748 1182 2751
rect 1202 2748 1214 2751
rect 1242 2748 1318 2751
rect 1322 2748 1430 2751
rect 1458 2748 1542 2751
rect 1546 2748 1734 2751
rect 1738 2748 1742 2751
rect 1850 2748 1862 2751
rect 1866 2748 2054 2751
rect 2066 2748 2118 2751
rect 2194 2748 2214 2751
rect 2222 2748 2230 2751
rect 2254 2751 2257 2758
rect 2254 2748 2281 2751
rect 2290 2748 2294 2751
rect 2414 2751 2417 2758
rect 2414 2748 2454 2751
rect 2482 2748 2510 2751
rect 2706 2748 2742 2751
rect 2746 2748 2982 2751
rect 3002 2748 3022 2751
rect 3182 2751 3185 2758
rect 3542 2752 3545 2758
rect 3146 2748 3185 2751
rect 3234 2748 3238 2751
rect 3258 2748 3286 2751
rect 3290 2748 3294 2751
rect 3314 2748 3409 2751
rect 3450 2748 3510 2751
rect 3590 2751 3594 2752
rect 3562 2748 3594 2751
rect 766 2742 769 2748
rect 886 2742 889 2748
rect 926 2742 929 2748
rect 2190 2742 2193 2748
rect 2222 2742 2225 2748
rect 2278 2742 2281 2748
rect 18 2738 38 2741
rect 154 2738 182 2741
rect 194 2738 206 2741
rect 226 2738 270 2741
rect 274 2738 414 2741
rect 418 2738 502 2741
rect 554 2738 614 2741
rect 618 2738 630 2741
rect 698 2738 758 2741
rect 786 2738 798 2741
rect 818 2738 838 2741
rect 874 2738 878 2741
rect 898 2738 918 2741
rect 974 2738 982 2741
rect 986 2738 1094 2741
rect 1178 2738 1302 2741
rect 1314 2738 1334 2741
rect 1514 2738 1566 2741
rect 1570 2738 1630 2741
rect 1634 2738 1662 2741
rect 1666 2738 1854 2741
rect 1858 2738 1910 2741
rect 1970 2738 1977 2741
rect 26 2728 54 2731
rect 138 2728 278 2731
rect 282 2728 358 2731
rect 482 2728 486 2731
rect 534 2728 537 2738
rect 694 2732 697 2738
rect 1422 2732 1425 2738
rect 1462 2732 1465 2738
rect 1974 2732 1977 2738
rect 2074 2738 2078 2741
rect 2082 2738 2110 2741
rect 2282 2738 2334 2741
rect 2342 2741 2345 2748
rect 2382 2741 2385 2748
rect 2638 2742 2641 2748
rect 2342 2738 2385 2741
rect 2426 2738 2462 2741
rect 2466 2738 2486 2741
rect 2506 2738 2574 2741
rect 2662 2741 2665 2748
rect 3406 2742 3409 2748
rect 2642 2738 2665 2741
rect 2802 2738 2814 2741
rect 2834 2738 2838 2741
rect 2850 2738 2862 2741
rect 2890 2738 2894 2741
rect 2994 2738 3086 2741
rect 3122 2738 3358 2741
rect 3386 2738 3398 2741
rect 3450 2738 3462 2741
rect 546 2728 566 2731
rect 650 2728 654 2731
rect 710 2728 718 2731
rect 722 2728 734 2731
rect 834 2728 1038 2731
rect 1106 2728 1110 2731
rect 1178 2728 1190 2731
rect 1298 2728 1326 2731
rect 1334 2728 1342 2731
rect 1346 2728 1358 2731
rect 1370 2728 1398 2731
rect 1578 2728 1582 2731
rect 1634 2728 1638 2731
rect 1658 2728 1710 2731
rect 1714 2728 1726 2731
rect 1738 2728 1806 2731
rect 1898 2728 1969 2731
rect 2038 2731 2041 2738
rect 2790 2732 2793 2738
rect 2038 2728 2078 2731
rect 2082 2728 2086 2731
rect 2114 2728 2118 2731
rect 2122 2728 2134 2731
rect 2186 2728 2198 2731
rect 2330 2728 2350 2731
rect 2802 2728 2822 2731
rect 2826 2728 2926 2731
rect 3034 2728 3054 2731
rect 3170 2728 3190 2731
rect 3202 2728 3230 2731
rect 3238 2728 3278 2731
rect 3282 2728 3318 2731
rect 3346 2728 3478 2731
rect 3590 2731 3594 2732
rect 3530 2728 3594 2731
rect 282 2718 286 2721
rect 354 2718 358 2721
rect 1054 2721 1057 2728
rect 370 2718 1057 2721
rect 1422 2721 1425 2728
rect 1066 2718 1425 2721
rect 1502 2721 1505 2728
rect 1502 2718 1574 2721
rect 1578 2718 1606 2721
rect 1610 2718 1646 2721
rect 1674 2718 1758 2721
rect 1778 2718 1798 2721
rect 1802 2718 1902 2721
rect 1906 2718 1926 2721
rect 1966 2721 1969 2728
rect 2006 2722 2009 2728
rect 2438 2722 2441 2728
rect 1966 2718 1990 2721
rect 2122 2718 2126 2721
rect 2226 2718 2318 2721
rect 2614 2721 2617 2728
rect 2530 2718 2617 2721
rect 2634 2718 2670 2721
rect 2766 2721 2769 2728
rect 2722 2718 2769 2721
rect 2794 2718 2934 2721
rect 2954 2718 2958 2721
rect 3034 2718 3038 2721
rect 3238 2721 3241 2728
rect 3202 2718 3241 2721
rect 3250 2718 3270 2721
rect 3290 2718 3294 2721
rect 3330 2718 3358 2721
rect 3450 2718 3518 2721
rect 194 2708 342 2711
rect 346 2708 446 2711
rect 474 2708 494 2711
rect 514 2708 550 2711
rect 554 2708 702 2711
rect 706 2708 726 2711
rect 762 2708 950 2711
rect 1050 2708 1086 2711
rect 1234 2708 1326 2711
rect 1338 2708 1350 2711
rect 1362 2708 1414 2711
rect 1418 2708 1446 2711
rect 1474 2708 1598 2711
rect 1618 2708 1630 2711
rect 1634 2708 1782 2711
rect 1794 2708 1974 2711
rect 2242 2708 2350 2711
rect 2434 2708 2590 2711
rect 2602 2708 2662 2711
rect 2714 2708 2742 2711
rect 2746 2708 2846 2711
rect 2938 2708 2950 2711
rect 2978 2708 3022 2711
rect 3326 2711 3329 2718
rect 3162 2708 3329 2711
rect 3410 2708 3486 2711
rect 3590 2711 3594 2712
rect 3490 2708 3594 2711
rect 992 2703 994 2707
rect 998 2703 1001 2707
rect 1006 2703 1008 2707
rect 2024 2703 2026 2707
rect 2030 2703 2033 2707
rect 2038 2703 2040 2707
rect 3040 2703 3042 2707
rect 3046 2703 3049 2707
rect 3054 2703 3056 2707
rect -26 2701 -22 2702
rect -26 2698 6 2701
rect 10 2698 30 2701
rect 34 2698 118 2701
rect 202 2698 270 2701
rect 274 2698 294 2701
rect 298 2698 318 2701
rect 330 2698 374 2701
rect 458 2698 510 2701
rect 522 2698 558 2701
rect 618 2698 654 2701
rect 666 2698 670 2701
rect 690 2698 718 2701
rect 842 2698 878 2701
rect 898 2698 902 2701
rect 922 2698 926 2701
rect 1042 2698 1142 2701
rect 1226 2698 1230 2701
rect 1258 2698 1918 2701
rect 1986 2698 2017 2701
rect 2226 2698 2342 2701
rect 2354 2698 2358 2701
rect 2554 2698 2598 2701
rect 2618 2698 2646 2701
rect 2658 2698 2830 2701
rect 2874 2698 2894 2701
rect 2914 2698 2982 2701
rect 3106 2698 3150 2701
rect 3154 2698 3174 2701
rect 3178 2698 3350 2701
rect 3354 2698 3494 2701
rect 10 2688 94 2691
rect 98 2688 214 2691
rect 374 2688 406 2691
rect 426 2688 446 2691
rect 450 2688 590 2691
rect 594 2688 902 2691
rect 926 2688 934 2691
rect 938 2688 1094 2691
rect 1114 2688 1262 2691
rect 1266 2688 1406 2691
rect 1474 2688 1534 2691
rect 1674 2688 1694 2691
rect 1834 2688 1838 2691
rect 1918 2688 1966 2691
rect 2002 2688 2006 2691
rect 2014 2691 2017 2698
rect 2014 2688 2254 2691
rect 2306 2688 2382 2691
rect 2402 2688 2638 2691
rect 2730 2688 2750 2691
rect 2758 2688 2766 2691
rect 2778 2688 2806 2691
rect 2818 2688 2838 2691
rect 2850 2688 2878 2691
rect 3034 2688 3038 2691
rect 3210 2688 3310 2691
rect 3318 2688 3366 2691
rect 3590 2691 3594 2692
rect 3562 2688 3594 2691
rect 374 2682 377 2688
rect 162 2678 206 2681
rect 234 2678 246 2681
rect 266 2678 374 2681
rect 394 2678 414 2681
rect 450 2678 454 2681
rect 466 2678 526 2681
rect 562 2678 566 2681
rect 578 2678 638 2681
rect 642 2678 694 2681
rect 746 2678 750 2681
rect 802 2678 1270 2681
rect 1386 2678 1414 2681
rect 1530 2678 1590 2681
rect 1658 2678 1670 2681
rect 1726 2681 1729 2688
rect 1686 2678 1729 2681
rect 1738 2678 1750 2681
rect 1754 2678 1782 2681
rect 1810 2678 1822 2681
rect 1898 2678 1910 2681
rect 1918 2681 1921 2688
rect 1914 2678 2062 2681
rect 2066 2678 2158 2681
rect 2170 2678 2206 2681
rect 2242 2678 2246 2681
rect 2346 2678 2350 2681
rect 2370 2678 2582 2681
rect 2586 2678 2678 2681
rect 2682 2678 2854 2681
rect 2874 2678 2910 2681
rect 2922 2678 2942 2681
rect 2986 2678 2990 2681
rect 3234 2678 3286 2681
rect 3318 2681 3321 2688
rect 3290 2678 3321 2681
rect 3378 2678 3390 2681
rect 3422 2681 3425 2688
rect 3394 2678 3425 2681
rect 3430 2681 3433 2688
rect 3478 2681 3481 2688
rect 3430 2678 3481 2681
rect 3498 2678 3593 2681
rect 14 2672 17 2678
rect 1686 2672 1689 2678
rect 26 2668 30 2671
rect 82 2668 150 2671
rect 170 2668 190 2671
rect 210 2668 286 2671
rect 338 2668 414 2671
rect 418 2668 942 2671
rect 946 2668 1134 2671
rect 1146 2668 1150 2671
rect 1162 2668 1166 2671
rect 1178 2668 1230 2671
rect 1274 2668 1422 2671
rect 1426 2668 1470 2671
rect 1570 2668 1598 2671
rect 1618 2668 1622 2671
rect 1650 2668 1678 2671
rect 1722 2668 1758 2671
rect 1762 2668 1886 2671
rect 1906 2668 1918 2671
rect 1922 2668 1942 2671
rect 1962 2668 1966 2671
rect 2106 2668 2118 2671
rect 2130 2668 2190 2671
rect 2310 2671 2313 2678
rect 3590 2672 3593 2678
rect 2226 2668 2313 2671
rect 2322 2668 2342 2671
rect 2402 2668 2406 2671
rect 2418 2670 2425 2671
rect 2418 2668 2422 2670
rect 18 2658 22 2661
rect 42 2658 54 2661
rect 66 2658 86 2661
rect 154 2658 230 2661
rect 234 2658 318 2661
rect 326 2661 329 2668
rect 2466 2668 2494 2671
rect 2506 2668 2534 2671
rect 2562 2668 2574 2671
rect 2594 2668 2625 2671
rect 2622 2662 2625 2668
rect 2642 2668 2689 2671
rect 2738 2668 2742 2671
rect 2762 2668 2766 2671
rect 2802 2668 2814 2671
rect 2826 2668 2830 2671
rect 2834 2668 2846 2671
rect 2874 2668 2998 2671
rect 3018 2668 3078 2671
rect 3202 2668 3262 2671
rect 3338 2668 3414 2671
rect 3418 2668 3446 2671
rect 3450 2668 3558 2671
rect 3590 2668 3594 2672
rect 2630 2662 2633 2668
rect 2686 2662 2689 2668
rect 326 2658 382 2661
rect 442 2658 510 2661
rect 530 2658 598 2661
rect 602 2658 622 2661
rect 650 2658 654 2661
rect 738 2658 750 2661
rect 762 2658 766 2661
rect 810 2658 830 2661
rect 834 2658 910 2661
rect 914 2658 934 2661
rect 954 2658 1038 2661
rect 1058 2658 1062 2661
rect 1114 2658 1126 2661
rect 1138 2658 1182 2661
rect 1218 2658 1246 2661
rect 1282 2658 1446 2661
rect 1458 2658 1486 2661
rect 1506 2658 1510 2661
rect 1698 2658 1734 2661
rect 1874 2658 2094 2661
rect 2106 2658 2118 2661
rect 2130 2658 2134 2661
rect 2138 2658 2150 2661
rect 2154 2658 2182 2661
rect 2186 2658 2518 2661
rect 2570 2658 2582 2661
rect 2586 2658 2606 2661
rect 2698 2658 2734 2661
rect 2782 2661 2785 2668
rect 3182 2662 3185 2668
rect 3270 2662 3273 2668
rect 3334 2662 3337 2668
rect 2778 2658 2785 2661
rect 2834 2658 2838 2661
rect 2858 2658 2862 2661
rect 2906 2658 2982 2661
rect 2994 2658 3134 2661
rect 3138 2658 3150 2661
rect 3394 2658 3417 2661
rect -26 2651 -22 2652
rect -26 2648 6 2651
rect 34 2648 78 2651
rect 122 2648 166 2651
rect 194 2648 222 2651
rect 298 2648 334 2651
rect 442 2648 446 2651
rect 538 2648 558 2651
rect 594 2648 598 2651
rect 770 2648 774 2651
rect 786 2648 1230 2651
rect 1322 2648 1409 2651
rect 1418 2648 1486 2651
rect 1534 2648 1542 2651
rect 1546 2648 1558 2651
rect 1574 2651 1577 2658
rect 1574 2648 1598 2651
rect 1626 2648 1638 2651
rect 1730 2648 1774 2651
rect 1778 2648 1854 2651
rect 1890 2648 1902 2651
rect 2026 2648 2054 2651
rect 2146 2648 2638 2651
rect 2642 2648 2710 2651
rect 2782 2651 2785 2658
rect 3414 2652 3417 2658
rect 2782 2648 2846 2651
rect 2986 2648 2998 2651
rect 3002 2648 3086 2651
rect 3138 2648 3254 2651
rect 3290 2648 3406 2651
rect 226 2638 382 2641
rect 478 2641 481 2648
rect 606 2642 609 2648
rect 410 2638 542 2641
rect 554 2638 582 2641
rect 650 2638 678 2641
rect 702 2641 705 2648
rect 702 2638 806 2641
rect 826 2638 838 2641
rect 858 2638 878 2641
rect 886 2638 918 2641
rect 954 2638 1014 2641
rect 1146 2638 1374 2641
rect 1406 2641 1409 2648
rect 1406 2638 1526 2641
rect 1586 2638 1646 2641
rect 1650 2638 1774 2641
rect 1778 2638 1886 2641
rect 1890 2638 2014 2641
rect 2066 2638 2158 2641
rect 2218 2638 2222 2641
rect 2386 2638 2470 2641
rect 2530 2638 2574 2641
rect 2578 2638 2585 2641
rect 2650 2638 2654 2641
rect 2722 2638 2742 2641
rect 2770 2638 2806 2641
rect 2842 2638 3118 2641
rect 3286 2641 3289 2648
rect 3154 2638 3289 2641
rect 3322 2638 3518 2641
rect -26 2631 -22 2632
rect -26 2628 22 2631
rect 26 2628 30 2631
rect 34 2628 102 2631
rect 106 2628 126 2631
rect 274 2628 462 2631
rect 594 2628 598 2631
rect 686 2631 689 2638
rect 886 2632 889 2638
rect 926 2632 929 2638
rect 686 2628 718 2631
rect 762 2628 790 2631
rect 794 2628 846 2631
rect 866 2628 870 2631
rect 882 2628 886 2631
rect 902 2628 910 2631
rect 978 2628 1054 2631
rect 1058 2628 1214 2631
rect 1234 2628 2790 2631
rect 2858 2628 2998 2631
rect 3290 2628 3342 2631
rect 18 2618 142 2621
rect 186 2618 310 2621
rect 354 2618 814 2621
rect 818 2618 982 2621
rect 986 2618 1102 2621
rect 1106 2618 1678 2621
rect 1682 2618 1830 2621
rect 1842 2618 1910 2621
rect 1922 2618 2350 2621
rect 2434 2618 2494 2621
rect 2522 2618 2654 2621
rect 2810 2618 2966 2621
rect 3238 2621 3241 2628
rect 3226 2618 3241 2621
rect 3338 2618 3382 2621
rect -26 2611 -22 2612
rect -26 2608 6 2611
rect 10 2608 30 2611
rect 98 2608 238 2611
rect 266 2608 422 2611
rect 522 2608 574 2611
rect 690 2608 766 2611
rect 770 2608 782 2611
rect 786 2608 878 2611
rect 1034 2608 1054 2611
rect 1082 2608 1318 2611
rect 1554 2608 1614 2611
rect 1658 2608 1790 2611
rect 1794 2608 1846 2611
rect 1882 2608 1998 2611
rect 2042 2608 2230 2611
rect 2306 2608 2510 2611
rect 2594 2608 2598 2611
rect 2658 2608 2894 2611
rect 2938 2608 2942 2611
rect 2970 2608 3217 2611
rect 3226 2608 3406 2611
rect 3410 2608 3438 2611
rect 480 2603 482 2607
rect 486 2603 489 2607
rect 494 2603 496 2607
rect 1512 2603 1514 2607
rect 1518 2603 1521 2607
rect 1526 2603 1528 2607
rect 2536 2603 2538 2607
rect 2542 2603 2545 2607
rect 2550 2603 2552 2607
rect 106 2598 358 2601
rect 562 2598 750 2601
rect 834 2598 846 2601
rect 882 2598 1174 2601
rect 1242 2598 1302 2601
rect 1314 2598 1454 2601
rect 1578 2598 1590 2601
rect 1682 2598 1710 2601
rect 1842 2598 1846 2601
rect 1866 2598 2006 2601
rect 2010 2598 2222 2601
rect 2410 2598 2526 2601
rect 2562 2598 2918 2601
rect 2938 2598 3206 2601
rect 3214 2601 3217 2608
rect 3214 2598 3374 2601
rect 3426 2598 3438 2601
rect -26 2591 -22 2592
rect -26 2588 142 2591
rect 174 2588 230 2591
rect 398 2591 401 2598
rect 438 2591 441 2598
rect 1478 2592 1481 2598
rect 398 2588 441 2591
rect 458 2588 534 2591
rect 618 2588 622 2591
rect 794 2588 958 2591
rect 962 2588 1086 2591
rect 1090 2588 1142 2591
rect 1186 2588 1286 2591
rect 1290 2588 1297 2591
rect 1338 2588 1430 2591
rect 1514 2588 1550 2591
rect 1562 2588 1798 2591
rect 1826 2588 1846 2591
rect 1874 2588 2854 2591
rect 2890 2588 3006 2591
rect 3042 2588 3142 2591
rect 3246 2588 3526 2591
rect 174 2582 177 2588
rect 218 2578 302 2581
rect 306 2578 334 2581
rect 362 2578 510 2581
rect 646 2581 649 2588
rect 3246 2582 3249 2588
rect 646 2578 830 2581
rect 834 2578 878 2581
rect 898 2578 902 2581
rect 914 2578 1310 2581
rect 1354 2578 1390 2581
rect 1410 2578 1758 2581
rect 1794 2578 1822 2581
rect 1826 2578 2054 2581
rect 2106 2578 2262 2581
rect 2330 2578 2558 2581
rect 2582 2578 2590 2581
rect 2594 2578 2606 2581
rect 2618 2578 2622 2581
rect 2698 2578 2814 2581
rect 2886 2578 2926 2581
rect 3082 2578 3110 2581
rect 3114 2578 3198 2581
rect 3346 2578 3462 2581
rect 3590 2581 3594 2582
rect 3562 2578 3594 2581
rect -26 2571 -22 2572
rect -26 2568 78 2571
rect 138 2568 190 2571
rect 330 2568 390 2571
rect 450 2568 566 2571
rect 586 2568 630 2571
rect 782 2568 1254 2571
rect 1306 2568 1390 2571
rect 1394 2568 1422 2571
rect 1426 2568 1897 2571
rect 2010 2568 2014 2571
rect 2154 2568 2174 2571
rect 2178 2568 2310 2571
rect 2434 2568 2438 2571
rect 2562 2568 2726 2571
rect 2886 2571 2889 2578
rect 2814 2568 2889 2571
rect 2958 2571 2961 2578
rect 2898 2568 2961 2571
rect 2978 2568 3014 2571
rect 3018 2568 3046 2571
rect 3202 2568 3350 2571
rect 3370 2568 3398 2571
rect 10 2558 62 2561
rect 126 2561 129 2568
rect 126 2558 238 2561
rect 242 2558 313 2561
rect 322 2558 326 2561
rect 514 2558 590 2561
rect 622 2558 718 2561
rect 726 2561 729 2568
rect 782 2562 785 2568
rect 1894 2562 1897 2568
rect 2814 2562 2817 2568
rect 726 2558 766 2561
rect 810 2558 838 2561
rect 842 2558 846 2561
rect 882 2558 1038 2561
rect 1074 2558 1086 2561
rect 1114 2558 1118 2561
rect 1178 2558 1190 2561
rect 1350 2558 1358 2561
rect 1362 2558 1454 2561
rect 1458 2558 1510 2561
rect 1530 2558 1646 2561
rect 1650 2558 1694 2561
rect 1706 2558 1761 2561
rect 1770 2558 1774 2561
rect 1826 2558 1886 2561
rect 1898 2558 2262 2561
rect 2290 2558 2334 2561
rect 2338 2558 2342 2561
rect 2458 2558 2462 2561
rect 2466 2558 2486 2561
rect 2506 2558 2526 2561
rect 2674 2558 2798 2561
rect 2922 2558 2950 2561
rect 2954 2558 3070 2561
rect 3106 2558 3182 2561
rect 3590 2561 3594 2562
rect 3426 2558 3594 2561
rect -26 2551 -22 2552
rect -26 2548 6 2551
rect 82 2548 134 2551
rect 282 2548 286 2551
rect 310 2551 313 2558
rect 430 2552 433 2558
rect 310 2548 382 2551
rect 474 2548 529 2551
rect 526 2542 529 2548
rect 614 2551 617 2558
rect 570 2548 617 2551
rect 622 2552 625 2558
rect 1214 2552 1217 2558
rect 1694 2552 1697 2558
rect 1758 2552 1761 2558
rect 2350 2552 2353 2558
rect 722 2548 734 2551
rect 738 2548 782 2551
rect 922 2548 942 2551
rect 946 2548 974 2551
rect 978 2548 1022 2551
rect 1026 2548 1118 2551
rect 1130 2548 1174 2551
rect 1322 2548 1366 2551
rect 1434 2548 1438 2551
rect 1442 2548 1454 2551
rect 1474 2548 1518 2551
rect 1538 2548 1558 2551
rect 1578 2548 1622 2551
rect 1674 2548 1678 2551
rect 1722 2548 1726 2551
rect 1738 2548 1742 2551
rect 1834 2548 1854 2551
rect 1930 2548 1958 2551
rect 2010 2548 2030 2551
rect 2034 2548 2046 2551
rect 2130 2548 2190 2551
rect 2226 2548 2278 2551
rect 2298 2548 2318 2551
rect 2322 2548 2350 2551
rect 2442 2548 2614 2551
rect 2618 2548 2734 2551
rect 2738 2548 2774 2551
rect 2874 2548 2878 2551
rect 3010 2548 3150 2551
rect 3290 2548 3318 2551
rect 3358 2548 3390 2551
rect 534 2542 537 2548
rect 10 2538 46 2541
rect 50 2538 166 2541
rect 170 2538 286 2541
rect 290 2538 350 2541
rect 354 2538 366 2541
rect 378 2538 470 2541
rect 490 2538 518 2541
rect 586 2538 614 2541
rect 618 2538 670 2541
rect 674 2538 710 2541
rect 722 2538 750 2541
rect 922 2538 934 2541
rect 946 2538 950 2541
rect 1002 2538 1006 2541
rect 1034 2538 1038 2541
rect 1074 2538 1078 2541
rect 1098 2540 1126 2541
rect 1094 2538 1126 2540
rect 1146 2538 1150 2541
rect 1178 2538 1318 2541
rect 1370 2538 1454 2541
rect 1554 2538 1566 2541
rect 1570 2538 1686 2541
rect 1690 2538 1734 2541
rect 1786 2538 1790 2541
rect 1834 2538 1838 2541
rect 1842 2538 1862 2541
rect 1890 2538 1894 2541
rect 1938 2538 1966 2541
rect 2050 2538 2070 2541
rect 2086 2538 2161 2541
rect 2170 2538 2209 2541
rect 34 2528 46 2531
rect 74 2528 278 2531
rect 290 2528 686 2531
rect 690 2528 702 2531
rect 746 2528 814 2531
rect 834 2528 862 2531
rect 898 2528 958 2531
rect 962 2528 998 2531
rect 1130 2528 1134 2531
rect 1282 2528 1406 2531
rect 1426 2528 1470 2531
rect 1522 2528 1606 2531
rect 1618 2528 1686 2531
rect 1910 2531 1913 2538
rect 1982 2532 1985 2538
rect 2086 2532 2089 2538
rect 2158 2532 2161 2538
rect 2206 2532 2209 2538
rect 2410 2538 2478 2541
rect 2490 2538 2494 2541
rect 2610 2538 2654 2541
rect 2690 2538 2710 2541
rect 2754 2538 2814 2541
rect 2842 2538 2846 2541
rect 2850 2538 3126 2541
rect 3154 2538 3158 2541
rect 3358 2541 3361 2548
rect 3162 2538 3361 2541
rect 3590 2541 3594 2542
rect 3378 2538 3594 2541
rect 2350 2532 2353 2538
rect 1690 2528 1918 2531
rect 2018 2528 2022 2531
rect 2066 2528 2070 2531
rect 2186 2528 2190 2531
rect 2210 2528 2214 2531
rect 2258 2528 2262 2531
rect 2410 2528 2470 2531
rect 2478 2531 2481 2538
rect 2590 2532 2593 2538
rect 2478 2528 2518 2531
rect 2530 2528 2534 2531
rect 2602 2528 2654 2531
rect 2658 2528 2750 2531
rect 3026 2528 3062 2531
rect 3146 2528 3174 2531
rect 3242 2528 3246 2531
rect 3266 2528 3342 2531
rect 1222 2522 1225 2528
rect 34 2518 62 2521
rect 74 2518 86 2521
rect 90 2518 110 2521
rect 154 2518 158 2521
rect 170 2518 222 2521
rect 318 2518 326 2521
rect 330 2518 334 2521
rect 370 2518 374 2521
rect 378 2518 406 2521
rect 434 2518 446 2521
rect 454 2518 462 2521
rect 466 2518 502 2521
rect 610 2518 614 2521
rect 682 2518 774 2521
rect 874 2518 1062 2521
rect 1102 2518 1110 2521
rect 1114 2518 1198 2521
rect 1362 2518 1454 2521
rect 1458 2518 1606 2521
rect 1610 2518 1654 2521
rect 1738 2518 1846 2521
rect 1858 2518 1926 2521
rect 1946 2518 2049 2521
rect 2058 2518 2174 2521
rect 2254 2521 2257 2528
rect 2398 2522 2401 2528
rect 2202 2518 2257 2521
rect 2290 2518 2382 2521
rect 2434 2518 2438 2521
rect 2458 2518 2478 2521
rect 2482 2518 2678 2521
rect 2730 2518 2838 2521
rect 3002 2518 3110 2521
rect 3146 2518 3182 2521
rect 3314 2518 3422 2521
rect 10 2508 142 2511
rect 154 2508 182 2511
rect 202 2508 270 2511
rect 274 2508 302 2511
rect 546 2508 574 2511
rect 586 2508 814 2511
rect 818 2508 846 2511
rect 850 2508 974 2511
rect 1034 2508 1086 2511
rect 1122 2508 1174 2511
rect 1290 2508 1334 2511
rect 1362 2508 1406 2511
rect 1482 2508 1558 2511
rect 1626 2508 1630 2511
rect 1650 2508 1718 2511
rect 1786 2508 1926 2511
rect 2046 2511 2049 2518
rect 2046 2508 2078 2511
rect 2162 2508 2374 2511
rect 2378 2508 2390 2511
rect 2402 2508 2414 2511
rect 2474 2508 2510 2511
rect 2514 2508 2566 2511
rect 2714 2508 2950 2511
rect 2954 2508 3014 2511
rect 3154 2508 3158 2511
rect 3170 2508 3286 2511
rect 992 2503 994 2507
rect 998 2503 1001 2507
rect 1006 2503 1008 2507
rect 2024 2503 2026 2507
rect 2030 2503 2033 2507
rect 2038 2503 2040 2507
rect 3040 2503 3042 2507
rect 3046 2503 3049 2507
rect 3054 2503 3056 2507
rect 42 2498 54 2501
rect 162 2498 198 2501
rect 210 2498 214 2501
rect 226 2498 262 2501
rect 266 2498 342 2501
rect 346 2498 454 2501
rect 466 2498 630 2501
rect 762 2498 798 2501
rect 802 2498 806 2501
rect 1018 2498 1062 2501
rect 1130 2498 1246 2501
rect 1330 2498 1334 2501
rect 1450 2498 1470 2501
rect 1474 2498 1502 2501
rect 1506 2498 1598 2501
rect 1602 2498 1654 2501
rect 1666 2498 1686 2501
rect 1738 2498 1790 2501
rect 1794 2498 1942 2501
rect 1946 2498 1990 2501
rect 2050 2498 2054 2501
rect 2062 2498 2070 2501
rect 2138 2498 2254 2501
rect 2466 2498 2510 2501
rect 2546 2498 2582 2501
rect 2586 2498 2598 2501
rect 2650 2498 2694 2501
rect 2698 2498 2734 2501
rect 2850 2498 2862 2501
rect 2866 2498 2934 2501
rect 3106 2498 3126 2501
rect 3130 2498 3310 2501
rect 1254 2492 1257 2498
rect 1374 2492 1377 2498
rect -26 2491 -22 2492
rect -26 2488 6 2491
rect 46 2488 86 2491
rect 90 2488 182 2491
rect 186 2488 206 2491
rect 410 2488 550 2491
rect 570 2488 598 2491
rect 714 2488 774 2491
rect 986 2488 1006 2491
rect 1058 2488 1062 2491
rect 1082 2488 1118 2491
rect 1170 2488 1246 2491
rect 1266 2488 1326 2491
rect 1446 2488 1454 2491
rect 1458 2488 1582 2491
rect 1594 2488 1630 2491
rect 1658 2488 1662 2491
rect 1754 2488 1766 2491
rect 1778 2488 1790 2491
rect 1826 2488 1830 2491
rect 1958 2488 1966 2491
rect 1970 2488 1990 2491
rect 2062 2491 2065 2498
rect 2010 2488 2065 2491
rect 2082 2488 2102 2491
rect 2154 2488 2209 2491
rect 2330 2488 2342 2491
rect 2458 2488 2526 2491
rect 2578 2488 2582 2491
rect 2594 2488 2598 2491
rect 2626 2488 2630 2491
rect 2730 2488 2886 2491
rect 2954 2488 3030 2491
rect 3122 2488 3126 2491
rect 3170 2488 3198 2491
rect 3286 2488 3294 2491
rect 3298 2488 3334 2491
rect 46 2482 49 2488
rect 606 2482 609 2488
rect 1406 2482 1409 2488
rect 1678 2482 1681 2488
rect 18 2478 30 2481
rect 58 2478 134 2481
rect 178 2478 198 2481
rect 322 2478 326 2481
rect 466 2478 470 2481
rect 498 2478 598 2481
rect 666 2478 686 2481
rect 698 2478 766 2481
rect 770 2478 1062 2481
rect 1106 2478 1206 2481
rect 1258 2478 1294 2481
rect 1298 2478 1406 2481
rect 1418 2478 1462 2481
rect 1538 2478 1574 2481
rect 1586 2478 1622 2481
rect 1706 2478 1830 2481
rect 2070 2481 2073 2488
rect 2206 2482 2209 2488
rect 1938 2478 2073 2481
rect 2090 2478 2102 2481
rect 2258 2478 2998 2481
rect 3114 2478 3334 2481
rect 3370 2478 3374 2481
rect 3386 2478 3422 2481
rect 18 2468 22 2471
rect 150 2471 153 2478
rect 446 2472 449 2478
rect 130 2468 190 2471
rect 298 2468 302 2471
rect 402 2468 438 2471
rect 530 2468 782 2471
rect 786 2468 806 2471
rect 914 2468 926 2471
rect 1010 2468 1038 2471
rect 1162 2468 1238 2471
rect 1246 2468 1302 2471
rect 1378 2468 1382 2471
rect 1394 2468 1430 2471
rect 1434 2468 1486 2471
rect 1498 2468 1502 2471
rect 1538 2468 1558 2471
rect 1562 2468 1606 2471
rect 1642 2468 1822 2471
rect 1826 2468 1878 2471
rect 1882 2468 1910 2471
rect 1954 2468 1974 2471
rect 1994 2468 2006 2471
rect 2026 2468 2062 2471
rect 2066 2468 2070 2471
rect 2234 2468 2254 2471
rect 2322 2468 2342 2471
rect 2370 2468 2406 2471
rect 2442 2468 2454 2471
rect 2482 2468 2486 2471
rect 2514 2468 2638 2471
rect 2758 2468 2814 2471
rect 2834 2468 2902 2471
rect 2970 2468 2990 2471
rect 3042 2468 3070 2471
rect 3074 2468 3081 2471
rect 3122 2468 3166 2471
rect 3178 2468 3222 2471
rect 3226 2468 3254 2471
rect 3346 2468 3390 2471
rect 878 2462 881 2468
rect 18 2458 22 2461
rect 146 2458 166 2461
rect 170 2458 206 2461
rect 290 2458 518 2461
rect 570 2458 574 2461
rect 626 2458 662 2461
rect 674 2458 678 2461
rect 690 2458 705 2461
rect 754 2458 758 2461
rect 794 2458 822 2461
rect 842 2458 870 2461
rect 898 2458 902 2461
rect 906 2458 918 2461
rect 934 2461 937 2468
rect 1246 2462 1249 2468
rect 2758 2462 2761 2468
rect 934 2458 998 2461
rect 1002 2458 1070 2461
rect 1082 2458 1134 2461
rect 1162 2458 1230 2461
rect 1242 2458 1246 2461
rect 1266 2458 1286 2461
rect 1298 2458 1398 2461
rect 1402 2458 1406 2461
rect 1418 2458 2254 2461
rect 2298 2458 2446 2461
rect 2450 2458 2478 2461
rect 2482 2458 2486 2461
rect 2514 2458 2518 2461
rect 2546 2458 2550 2461
rect 2578 2458 2590 2461
rect 2626 2458 2718 2461
rect 2786 2458 2894 2461
rect 2954 2458 2958 2461
rect 3034 2458 3118 2461
rect 3126 2458 3142 2461
rect 3250 2458 3254 2461
rect 3418 2458 3422 2461
rect 3514 2458 3518 2461
rect -26 2451 -22 2452
rect -26 2448 54 2451
rect 66 2448 97 2451
rect 122 2448 150 2451
rect 318 2448 425 2451
rect 482 2448 502 2451
rect 546 2448 566 2451
rect 594 2448 694 2451
rect 702 2451 705 2458
rect 702 2448 766 2451
rect 818 2448 886 2451
rect 934 2451 937 2458
rect 2670 2452 2673 2458
rect 930 2448 937 2451
rect 954 2448 974 2451
rect 1058 2448 1094 2451
rect 1114 2448 1118 2451
rect 1122 2448 1214 2451
rect 1222 2448 1230 2451
rect 1234 2448 1286 2451
rect 1298 2448 1382 2451
rect 1386 2448 1438 2451
rect 1466 2448 1502 2451
rect 1522 2448 1526 2451
rect 1546 2448 1566 2451
rect 1586 2448 1590 2451
rect 1678 2448 1718 2451
rect 1738 2448 1742 2451
rect 1770 2448 1798 2451
rect 1814 2448 1822 2451
rect 1826 2448 2134 2451
rect 2194 2448 2222 2451
rect 2242 2448 2270 2451
rect 2290 2448 2297 2451
rect 2330 2448 2358 2451
rect 2370 2448 2470 2451
rect 2482 2448 2590 2451
rect 2730 2448 2766 2451
rect 2786 2448 2806 2451
rect 2818 2448 2854 2451
rect 2922 2448 2950 2451
rect 2962 2448 2969 2451
rect 3126 2451 3129 2458
rect 2986 2448 3129 2451
rect 3138 2448 3142 2451
rect 3194 2448 3198 2451
rect 3202 2448 3270 2451
rect 3274 2448 3342 2451
rect 3346 2448 3350 2451
rect 3354 2448 3366 2451
rect 3394 2448 3470 2451
rect 94 2442 97 2448
rect 318 2442 321 2448
rect 422 2442 425 2448
rect 138 2438 158 2441
rect 162 2438 230 2441
rect 234 2438 238 2441
rect 538 2438 758 2441
rect 770 2438 838 2441
rect 842 2438 870 2441
rect 886 2441 889 2448
rect 1678 2442 1681 2448
rect 2294 2442 2297 2448
rect 2966 2442 2969 2448
rect 3534 2442 3537 2448
rect 886 2438 966 2441
rect 978 2438 998 2441
rect 1002 2438 1014 2441
rect 1042 2438 1134 2441
rect 1186 2438 1190 2441
rect 1210 2438 1318 2441
rect 1322 2438 1326 2441
rect 1394 2438 1398 2441
rect 1522 2438 1550 2441
rect 1766 2438 1774 2441
rect 1778 2438 2086 2441
rect 2106 2438 2134 2441
rect 2138 2438 2158 2441
rect 2186 2438 2238 2441
rect 2254 2438 2262 2441
rect 2266 2438 2286 2441
rect 2342 2438 2350 2441
rect 2354 2438 2374 2441
rect 2522 2438 2542 2441
rect 2602 2438 2702 2441
rect 2706 2438 2742 2441
rect 2778 2438 2790 2441
rect 2842 2438 2870 2441
rect 3034 2438 3062 2441
rect 3146 2438 3302 2441
rect 66 2428 110 2431
rect 114 2428 134 2431
rect 138 2428 158 2431
rect 258 2428 414 2431
rect 418 2428 422 2431
rect 1142 2431 1145 2438
rect 514 2428 1145 2431
rect 1422 2431 1425 2438
rect 1186 2428 2414 2431
rect 2418 2428 2438 2431
rect 2530 2428 3118 2431
rect 3122 2428 3158 2431
rect 3186 2428 3230 2431
rect 3234 2428 3270 2431
rect 3274 2428 3278 2431
rect 146 2418 374 2421
rect 486 2421 489 2428
rect 458 2418 489 2421
rect 506 2418 678 2421
rect 698 2418 854 2421
rect 858 2418 865 2421
rect 970 2418 1574 2421
rect 1650 2418 1750 2421
rect 1810 2418 1838 2421
rect 1842 2418 1862 2421
rect 1890 2418 1958 2421
rect 1986 2418 2246 2421
rect 2250 2418 2574 2421
rect 2746 2418 2774 2421
rect 2890 2418 2894 2421
rect 2922 2418 3454 2421
rect 354 2408 470 2411
rect 850 2408 990 2411
rect 994 2408 1014 2411
rect 1074 2408 1166 2411
rect 1186 2408 1198 2411
rect 1234 2408 1273 2411
rect 1306 2408 1366 2411
rect 1370 2408 1398 2411
rect 1418 2408 1422 2411
rect 1554 2408 1702 2411
rect 1890 2408 1902 2411
rect 2074 2408 2198 2411
rect 2218 2408 2318 2411
rect 2378 2408 2390 2411
rect 2642 2408 2974 2411
rect 3058 2408 3094 2411
rect 480 2403 482 2407
rect 486 2403 489 2407
rect 494 2403 496 2407
rect -26 2401 -22 2402
rect -26 2398 6 2401
rect 314 2398 462 2401
rect 506 2398 558 2401
rect 586 2398 686 2401
rect 714 2398 758 2401
rect 970 2398 982 2401
rect 1026 2398 1030 2401
rect 1050 2398 1054 2401
rect 1130 2398 1214 2401
rect 1250 2398 1262 2401
rect 1270 2401 1273 2408
rect 1512 2403 1514 2407
rect 1518 2403 1521 2407
rect 1526 2403 1528 2407
rect 2536 2403 2538 2407
rect 2542 2403 2545 2407
rect 2550 2403 2552 2407
rect 1270 2398 1326 2401
rect 1378 2398 1390 2401
rect 1650 2398 2046 2401
rect 2154 2398 2382 2401
rect 2650 2398 2830 2401
rect 2858 2398 3102 2401
rect 3106 2398 3366 2401
rect 402 2388 438 2391
rect 466 2388 694 2391
rect 730 2388 878 2391
rect 918 2388 1462 2391
rect 1466 2388 1510 2391
rect 1514 2388 1542 2391
rect 1562 2388 1646 2391
rect 1658 2388 1686 2391
rect 1930 2388 2198 2391
rect 2202 2388 2326 2391
rect 2394 2388 2398 2391
rect 2418 2388 2718 2391
rect 3094 2388 3134 2391
rect 918 2382 921 2388
rect 3094 2382 3097 2388
rect 34 2378 94 2381
rect 242 2378 321 2381
rect 318 2372 321 2378
rect 442 2378 518 2381
rect 586 2378 638 2381
rect 754 2378 766 2381
rect 794 2378 825 2381
rect 858 2378 886 2381
rect 1146 2378 1150 2381
rect 1170 2378 1278 2381
rect 1378 2378 1430 2381
rect 1434 2378 2854 2381
rect -26 2371 -22 2372
rect -26 2368 6 2371
rect 42 2368 54 2371
rect 122 2368 174 2371
rect 290 2368 294 2371
rect 342 2371 345 2378
rect 338 2368 345 2371
rect 354 2368 358 2371
rect 378 2368 582 2371
rect 706 2368 734 2371
rect 778 2368 814 2371
rect 822 2371 825 2378
rect 822 2368 910 2371
rect 1074 2368 1110 2371
rect 1122 2368 1134 2371
rect 1146 2368 1158 2371
rect 1194 2368 1214 2371
rect 1218 2368 1294 2371
rect 1346 2368 1446 2371
rect 1482 2368 1574 2371
rect 1778 2368 1878 2371
rect 1890 2368 1894 2371
rect 1914 2368 2054 2371
rect 2074 2368 2094 2371
rect 2230 2368 2238 2371
rect 2242 2368 2270 2371
rect 2282 2368 2366 2371
rect 2370 2368 2614 2371
rect 2618 2368 2686 2371
rect 2690 2368 2766 2371
rect 2786 2368 2830 2371
rect 2934 2371 2937 2378
rect 2874 2368 2937 2371
rect 3146 2368 3246 2371
rect 3294 2368 3334 2371
rect 62 2361 65 2368
rect 50 2358 65 2361
rect 106 2358 110 2361
rect 130 2358 214 2361
rect 218 2358 614 2361
rect 622 2358 630 2361
rect 638 2361 641 2368
rect 758 2362 761 2368
rect 2950 2362 2953 2368
rect 3294 2362 3297 2368
rect 638 2358 662 2361
rect 722 2358 726 2361
rect 826 2358 830 2361
rect 882 2358 902 2361
rect 954 2358 1022 2361
rect 1042 2358 1286 2361
rect 1290 2358 1398 2361
rect 1530 2358 1582 2361
rect 1610 2358 1614 2361
rect 1722 2358 1742 2361
rect 1802 2358 1974 2361
rect 2130 2358 2158 2361
rect 2194 2358 2470 2361
rect 2514 2358 2534 2361
rect 2538 2358 2582 2361
rect 2594 2358 2598 2361
rect 2610 2358 2630 2361
rect 2658 2358 2742 2361
rect 2826 2358 2918 2361
rect 2922 2358 2942 2361
rect 2970 2358 2974 2361
rect 3202 2358 3214 2361
rect 3242 2358 3254 2361
rect 3330 2358 3350 2361
rect 3362 2358 3382 2361
rect 3402 2358 3406 2361
rect 3438 2361 3441 2368
rect 3438 2358 3462 2361
rect 622 2352 625 2358
rect -26 2351 -22 2352
rect -26 2348 6 2351
rect 34 2348 510 2351
rect 546 2348 550 2351
rect 682 2348 702 2351
rect 714 2348 782 2351
rect 794 2348 798 2351
rect 802 2348 862 2351
rect 866 2348 886 2351
rect 898 2348 910 2351
rect 914 2348 918 2351
rect 942 2351 945 2358
rect 1662 2352 1665 2358
rect 2110 2352 2113 2358
rect 938 2348 945 2351
rect 1010 2348 1046 2351
rect 1066 2348 1110 2351
rect 1114 2348 1230 2351
rect 1234 2348 1246 2351
rect 1274 2348 1302 2351
rect 1354 2348 1358 2351
rect 1418 2348 1454 2351
rect 1458 2348 1574 2351
rect 1650 2348 1654 2351
rect 1706 2348 1822 2351
rect 1826 2348 1894 2351
rect 1898 2348 1934 2351
rect 1978 2348 1982 2351
rect 1986 2348 1998 2351
rect 2002 2348 2030 2351
rect 2050 2348 2094 2351
rect 2202 2348 2222 2351
rect 2234 2348 2294 2351
rect 2298 2348 2310 2351
rect 2330 2348 2334 2351
rect 2386 2348 2422 2351
rect 2426 2348 2486 2351
rect 2594 2348 2654 2351
rect 2682 2348 2702 2351
rect 2746 2348 2870 2351
rect 2914 2348 2942 2351
rect 2946 2348 2950 2351
rect 3042 2348 3086 2351
rect 3170 2348 3190 2351
rect 3210 2348 3334 2351
rect 3338 2348 3494 2351
rect 3498 2348 3502 2351
rect 3590 2351 3594 2352
rect 3562 2348 3594 2351
rect 654 2342 657 2348
rect 1254 2342 1257 2348
rect 1334 2342 1337 2348
rect 1406 2342 1409 2348
rect 34 2338 38 2341
rect 106 2338 390 2341
rect 394 2338 398 2341
rect 410 2338 414 2341
rect 426 2338 438 2341
rect 442 2338 470 2341
rect 514 2338 534 2341
rect 538 2338 542 2341
rect 562 2338 598 2341
rect 602 2338 654 2341
rect 666 2338 670 2341
rect 690 2338 766 2341
rect 786 2338 790 2341
rect 818 2338 822 2341
rect 834 2338 918 2341
rect 922 2338 974 2341
rect 978 2338 1094 2341
rect 1098 2338 1134 2341
rect 1138 2338 1142 2341
rect 1170 2338 1198 2341
rect 1218 2338 1246 2341
rect 1498 2338 1502 2341
rect 1610 2338 1718 2341
rect 1730 2338 1734 2341
rect 1746 2338 1750 2341
rect 1754 2338 1766 2341
rect 1778 2338 1782 2341
rect 1802 2338 1918 2341
rect 1922 2338 1942 2341
rect 2002 2338 2166 2341
rect 2170 2338 2225 2341
rect 2266 2338 2270 2341
rect 2274 2338 2350 2341
rect 2402 2338 2654 2341
rect 2658 2338 2774 2341
rect 2778 2338 2862 2341
rect 2930 2338 2934 2341
rect 2946 2338 3094 2341
rect 3122 2338 3126 2341
rect 3170 2338 3198 2341
rect 3202 2338 3238 2341
rect 3242 2338 3318 2341
rect 3386 2338 3390 2341
rect 3418 2338 3430 2341
rect 3466 2338 3478 2341
rect 82 2328 174 2331
rect 186 2328 190 2331
rect 306 2328 334 2331
rect 346 2328 350 2331
rect 370 2328 374 2331
rect 386 2328 414 2331
rect 434 2328 486 2331
rect 530 2328 534 2331
rect 830 2331 833 2338
rect 1950 2332 1953 2338
rect 2222 2332 2225 2338
rect 3366 2332 3369 2338
rect 3446 2332 3449 2338
rect 618 2328 833 2331
rect 874 2328 1046 2331
rect 1050 2328 1134 2331
rect 1170 2328 1358 2331
rect 1522 2328 1526 2331
rect 1642 2328 1710 2331
rect 1746 2328 1758 2331
rect 1778 2328 1782 2331
rect 1842 2328 1846 2331
rect 1874 2328 1902 2331
rect 2010 2328 2070 2331
rect 2090 2328 2094 2331
rect 2098 2328 2102 2331
rect 2114 2328 2134 2331
rect 2362 2328 2446 2331
rect 2474 2328 2494 2331
rect 2506 2328 2510 2331
rect 2562 2328 2566 2331
rect 2586 2328 2598 2331
rect 2650 2328 2670 2331
rect 2754 2328 2806 2331
rect 2842 2328 2862 2331
rect 2890 2328 2950 2331
rect 3018 2328 3230 2331
rect 3322 2328 3326 2331
rect 3338 2328 3350 2331
rect 3386 2328 3446 2331
rect 178 2318 198 2321
rect 202 2318 222 2321
rect 234 2318 406 2321
rect 410 2318 550 2321
rect 570 2318 574 2321
rect 602 2318 646 2321
rect 654 2318 710 2321
rect 722 2318 726 2321
rect 738 2318 742 2321
rect 758 2318 766 2321
rect 770 2318 782 2321
rect 854 2321 857 2328
rect 810 2318 857 2321
rect 866 2318 870 2321
rect 878 2318 1326 2321
rect 1330 2318 2006 2321
rect 2018 2318 2142 2321
rect 2262 2321 2265 2328
rect 2694 2322 2697 2328
rect 2146 2318 2265 2321
rect 2298 2318 2374 2321
rect 2490 2318 2550 2321
rect 2570 2318 2678 2321
rect 2862 2318 2870 2321
rect 2874 2318 2966 2321
rect 2978 2318 3054 2321
rect 3274 2318 3278 2321
rect 3314 2318 3414 2321
rect 154 2308 350 2311
rect 426 2308 438 2311
rect 498 2308 606 2311
rect 654 2311 657 2318
rect 618 2308 657 2311
rect 682 2308 694 2311
rect 878 2311 881 2318
rect 698 2308 881 2311
rect 962 2308 966 2311
rect 1018 2308 1150 2311
rect 1158 2308 1206 2311
rect 1218 2308 1222 2311
rect 1290 2308 1454 2311
rect 1594 2308 1790 2311
rect 1834 2308 1838 2311
rect 1946 2308 1998 2311
rect 2082 2308 2182 2311
rect 2418 2308 2726 2311
rect 2730 2308 2758 2311
rect 2766 2308 2822 2311
rect 2858 2308 2878 2311
rect 2906 2308 2918 2311
rect 3170 2308 3246 2311
rect 3258 2308 3334 2311
rect 3338 2308 3382 2311
rect 3394 2308 3422 2311
rect 3426 2308 3454 2311
rect 992 2303 994 2307
rect 998 2303 1001 2307
rect 1006 2303 1008 2307
rect 66 2298 102 2301
rect 226 2298 494 2301
rect 554 2298 558 2301
rect 634 2298 926 2301
rect 930 2298 982 2301
rect 1018 2298 1054 2301
rect 1158 2301 1161 2308
rect 1146 2298 1161 2301
rect 1178 2298 1222 2301
rect 1242 2298 1278 2301
rect 1290 2298 1342 2301
rect 1454 2301 1457 2308
rect 1454 2298 1598 2301
rect 1602 2298 1654 2301
rect 1658 2298 1726 2301
rect 1730 2298 1750 2301
rect 1762 2298 1766 2301
rect 1942 2301 1945 2308
rect 2024 2303 2026 2307
rect 2030 2303 2033 2307
rect 2038 2303 2040 2307
rect 1834 2298 1945 2301
rect 2050 2298 2222 2301
rect 2226 2298 2246 2301
rect 2250 2298 2254 2301
rect 2458 2298 2582 2301
rect 2594 2298 2638 2301
rect 2650 2298 2670 2301
rect 2766 2301 2769 2308
rect 3040 2303 3042 2307
rect 3046 2303 3049 2307
rect 3054 2303 3056 2307
rect 2682 2298 2769 2301
rect 2786 2298 2918 2301
rect 2938 2298 2982 2301
rect 2986 2298 2998 2301
rect 3178 2298 3414 2301
rect 3530 2298 3550 2301
rect 3590 2301 3594 2302
rect 3562 2298 3594 2301
rect 3134 2292 3137 2298
rect 130 2288 150 2291
rect 458 2288 542 2291
rect 546 2288 822 2291
rect 826 2288 934 2291
rect 938 2288 998 2291
rect 1002 2288 1118 2291
rect 1154 2288 1174 2291
rect 1178 2288 1238 2291
rect 1266 2288 1278 2291
rect 1402 2288 1430 2291
rect 1442 2288 1542 2291
rect 1570 2288 1630 2291
rect 1838 2288 1846 2291
rect 1850 2288 1894 2291
rect 1902 2288 1958 2291
rect 2014 2288 2158 2291
rect 2162 2288 2198 2291
rect 2442 2288 2622 2291
rect 2690 2288 2710 2291
rect 2714 2288 2854 2291
rect 2918 2288 2926 2291
rect 2930 2288 3102 2291
rect 3202 2288 3206 2291
rect 3218 2288 3318 2291
rect 3330 2288 3350 2291
rect 3370 2288 3374 2291
rect 3378 2288 3422 2291
rect 106 2278 246 2281
rect 282 2278 334 2281
rect 394 2278 574 2281
rect 602 2278 606 2281
rect 666 2278 718 2281
rect 762 2278 798 2281
rect 850 2278 902 2281
rect 954 2278 958 2281
rect 1042 2278 1046 2281
rect 1058 2278 1062 2281
rect 1106 2278 1118 2281
rect 1138 2278 1166 2281
rect 1186 2278 1190 2281
rect 1226 2278 1230 2281
rect 1274 2278 1278 2281
rect 1298 2278 1350 2281
rect 1450 2278 1454 2281
rect 1506 2278 1550 2281
rect 1554 2278 1566 2281
rect 1578 2278 1686 2281
rect 1722 2278 1726 2281
rect 1746 2278 1782 2281
rect 1786 2278 1798 2281
rect 1814 2281 1817 2288
rect 1902 2282 1905 2288
rect 2014 2282 2017 2288
rect 2326 2282 2329 2288
rect 1814 2278 1838 2281
rect 1962 2278 1966 2281
rect 1978 2278 2014 2281
rect 2146 2278 2150 2281
rect 2186 2278 2214 2281
rect 2382 2281 2385 2288
rect 2382 2278 2406 2281
rect 2410 2278 2422 2281
rect 2426 2278 2430 2281
rect 2458 2278 2462 2281
rect 2466 2278 2502 2281
rect 2578 2278 2582 2281
rect 2602 2278 2606 2281
rect 2666 2278 2702 2281
rect 2738 2278 2758 2281
rect 2762 2278 2766 2281
rect 2810 2278 2814 2281
rect 2914 2278 2998 2281
rect 3002 2278 3150 2281
rect 3162 2278 3214 2281
rect 3590 2281 3594 2282
rect 3218 2278 3594 2281
rect -26 2271 -22 2272
rect -26 2268 6 2271
rect 58 2268 78 2271
rect 98 2268 102 2271
rect 122 2268 134 2271
rect 186 2268 342 2271
rect 362 2268 366 2271
rect 434 2268 446 2271
rect 506 2268 518 2271
rect 554 2268 582 2271
rect 618 2268 686 2271
rect 762 2268 766 2271
rect 850 2268 854 2271
rect 882 2268 886 2271
rect 898 2268 918 2271
rect 922 2268 1062 2271
rect 1066 2268 1190 2271
rect 1194 2268 1246 2271
rect 1262 2271 1265 2278
rect 1262 2268 1294 2271
rect 1314 2268 1382 2271
rect 1430 2271 1433 2278
rect 1430 2268 1446 2271
rect 1474 2268 1534 2271
rect 1546 2268 1558 2271
rect 1578 2268 1582 2271
rect 1618 2268 1622 2271
rect 1658 2268 1694 2271
rect 1698 2268 1862 2271
rect 1878 2271 1881 2278
rect 2110 2272 2113 2278
rect 2126 2272 2129 2278
rect 1878 2268 1902 2271
rect 1906 2268 2014 2271
rect 2074 2268 2078 2271
rect 2138 2268 2166 2271
rect 2194 2268 2198 2271
rect 2210 2268 2214 2271
rect 2226 2270 2273 2271
rect 2226 2268 2270 2270
rect 2282 2268 2310 2271
rect 2314 2268 2318 2271
rect 2386 2268 2430 2271
rect 2434 2268 2478 2271
rect 2490 2268 2574 2271
rect 2642 2268 2742 2271
rect 2762 2268 3062 2271
rect 3066 2268 3126 2271
rect 3130 2268 3190 2271
rect 3210 2268 3310 2271
rect 3314 2268 3398 2271
rect 3402 2268 3454 2271
rect 3458 2268 3558 2271
rect 26 2258 38 2261
rect 42 2258 614 2261
rect 714 2258 806 2261
rect 810 2258 910 2261
rect 914 2258 1086 2261
rect 1090 2258 1094 2261
rect 1146 2258 1398 2261
rect 1458 2258 1606 2261
rect 1610 2258 1910 2261
rect 1946 2258 2022 2261
rect 2034 2258 2286 2261
rect 2290 2258 2390 2261
rect 2442 2258 2678 2261
rect 2706 2258 2713 2261
rect 2722 2258 2750 2261
rect 2770 2258 3054 2261
rect 3058 2258 3118 2261
rect 3122 2258 3158 2261
rect 3590 2261 3594 2262
rect 3194 2258 3594 2261
rect -26 2251 -22 2252
rect -26 2248 14 2251
rect 34 2248 94 2251
rect 138 2248 182 2251
rect 186 2248 230 2251
rect 234 2248 254 2251
rect 258 2248 302 2251
rect 306 2248 342 2251
rect 466 2248 526 2251
rect 570 2248 574 2251
rect 586 2248 646 2251
rect 690 2248 734 2251
rect 746 2248 750 2251
rect 754 2248 1142 2251
rect 1146 2248 1158 2251
rect 1162 2248 1166 2251
rect 1206 2248 1294 2251
rect 1338 2248 1374 2251
rect 1378 2248 1414 2251
rect 1442 2248 1470 2251
rect 1558 2248 1598 2251
rect 1602 2248 1686 2251
rect 1698 2248 1702 2251
rect 1714 2248 1750 2251
rect 1802 2248 1822 2251
rect 1970 2248 2238 2251
rect 2258 2248 2297 2251
rect 2306 2248 2310 2251
rect 2370 2248 2406 2251
rect 2426 2248 2446 2251
rect 2450 2248 2518 2251
rect 2610 2248 2638 2251
rect 2706 2248 2734 2251
rect 2770 2248 2854 2251
rect 2866 2248 2870 2251
rect 2906 2248 2950 2251
rect 3042 2248 3070 2251
rect 3090 2248 3094 2251
rect 3138 2248 3153 2251
rect 3178 2248 3214 2251
rect 3242 2248 3398 2251
rect 3402 2248 3446 2251
rect 3514 2248 3542 2251
rect 1206 2242 1209 2248
rect 1558 2242 1561 2248
rect 42 2238 54 2241
rect 338 2238 390 2241
rect 394 2238 510 2241
rect 530 2238 590 2241
rect 642 2238 662 2241
rect 682 2238 694 2241
rect 762 2238 870 2241
rect 874 2238 1006 2241
rect 1122 2238 1150 2241
rect 1250 2238 1278 2241
rect 1282 2238 1438 2241
rect 2294 2241 2297 2248
rect 3150 2242 3153 2248
rect 1642 2238 2281 2241
rect 2294 2238 2342 2241
rect 2498 2238 2502 2241
rect 2570 2238 2638 2241
rect 2746 2238 2886 2241
rect 2890 2238 3078 2241
rect 3154 2238 3182 2241
rect 3222 2241 3225 2248
rect 3210 2238 3225 2241
rect 3242 2238 3246 2241
rect 3290 2238 3318 2241
rect 3322 2238 3470 2241
rect 10 2228 782 2231
rect 786 2228 974 2231
rect 978 2228 1134 2231
rect 1138 2228 1174 2231
rect 1218 2228 1257 2231
rect 1354 2228 1502 2231
rect 1586 2228 2166 2231
rect 2178 2228 2270 2231
rect 2278 2231 2281 2238
rect 3286 2231 3289 2238
rect 2278 2228 3289 2231
rect 3298 2228 3342 2231
rect 3346 2228 3425 2231
rect 154 2218 502 2221
rect 562 2218 758 2221
rect 762 2218 1110 2221
rect 1190 2221 1193 2228
rect 1130 2218 1193 2221
rect 1254 2222 1257 2228
rect 3422 2222 3425 2228
rect 1446 2218 1654 2221
rect 1682 2218 2758 2221
rect 2762 2218 2806 2221
rect 2842 2218 2974 2221
rect 2978 2218 2990 2221
rect 3002 2218 3102 2221
rect 3106 2218 3174 2221
rect 3186 2218 3190 2221
rect 3242 2218 3246 2221
rect 3266 2218 3342 2221
rect 3346 2218 3390 2221
rect 170 2208 286 2211
rect 362 2208 446 2211
rect 594 2208 726 2211
rect 730 2208 1102 2211
rect 1446 2211 1449 2218
rect 1106 2208 1449 2211
rect 1714 2208 2062 2211
rect 2066 2208 2110 2211
rect 2114 2208 2118 2211
rect 2122 2208 2334 2211
rect 2514 2208 2518 2211
rect 2770 2208 2774 2211
rect 2802 2208 2918 2211
rect 2922 2208 2998 2211
rect 3226 2208 3422 2211
rect 480 2203 482 2207
rect 486 2203 489 2207
rect 494 2203 496 2207
rect 1512 2203 1514 2207
rect 1518 2203 1521 2207
rect 1526 2203 1528 2207
rect 2536 2203 2538 2207
rect 2542 2203 2545 2207
rect 2550 2203 2552 2207
rect 82 2198 238 2201
rect 274 2198 366 2201
rect 506 2198 582 2201
rect 658 2198 718 2201
rect 730 2198 798 2201
rect 818 2198 886 2201
rect 898 2198 958 2201
rect 962 2198 1078 2201
rect 1090 2198 1126 2201
rect 1170 2198 1265 2201
rect 1282 2198 1374 2201
rect 1458 2198 1486 2201
rect 1546 2198 1782 2201
rect 1794 2198 1798 2201
rect 1810 2198 1838 2201
rect 1882 2198 1886 2201
rect 1914 2198 1966 2201
rect 2018 2198 2062 2201
rect 2074 2198 2078 2201
rect 2090 2198 2198 2201
rect 2210 2198 2430 2201
rect 2570 2198 2798 2201
rect 2818 2198 2862 2201
rect 2954 2198 3430 2201
rect 3434 2198 3478 2201
rect 3590 2201 3594 2202
rect 3482 2198 3594 2201
rect 570 2188 918 2191
rect 962 2188 1230 2191
rect 1262 2191 1265 2198
rect 1262 2188 1310 2191
rect 1314 2188 1342 2191
rect 1378 2188 1718 2191
rect 1754 2188 2902 2191
rect 2938 2188 2977 2191
rect 3170 2188 3438 2191
rect 1718 2182 1721 2188
rect 2974 2182 2977 2188
rect -26 2181 -22 2182
rect -26 2178 81 2181
rect 114 2178 134 2181
rect 218 2178 342 2181
rect 346 2178 1382 2181
rect 1426 2178 1510 2181
rect 1538 2178 1542 2181
rect 1554 2178 1558 2181
rect 1618 2178 1670 2181
rect 1722 2178 1790 2181
rect 1794 2178 1830 2181
rect 1834 2178 1902 2181
rect 1914 2178 2270 2181
rect 2274 2178 2718 2181
rect 3026 2178 3110 2181
rect 3194 2178 3326 2181
rect 18 2168 22 2171
rect 78 2171 81 2178
rect 78 2168 190 2171
rect 282 2168 294 2171
rect 314 2168 318 2171
rect 370 2168 374 2171
rect 434 2168 478 2171
rect 482 2168 550 2171
rect 634 2168 638 2171
rect 682 2168 686 2171
rect 706 2168 822 2171
rect 858 2168 862 2171
rect 898 2168 902 2171
rect 946 2168 950 2171
rect 954 2168 982 2171
rect 994 2168 1014 2171
rect 1058 2168 1070 2171
rect 1098 2168 1166 2171
rect 1170 2168 1662 2171
rect 1666 2168 1886 2171
rect 1890 2168 1950 2171
rect 1954 2168 2030 2171
rect 2050 2168 2054 2171
rect 2106 2168 2134 2171
rect 2146 2168 2238 2171
rect 2386 2168 2406 2171
rect 2426 2168 2518 2171
rect 2546 2168 2654 2171
rect 2690 2168 2806 2171
rect 3242 2168 3310 2171
rect 3590 2171 3594 2172
rect 3458 2168 3594 2171
rect 2086 2162 2089 2168
rect -26 2161 -22 2162
rect -26 2158 30 2161
rect 34 2158 110 2161
rect 202 2158 278 2161
rect 314 2158 502 2161
rect 546 2158 550 2161
rect 586 2158 590 2161
rect 594 2158 790 2161
rect 794 2158 950 2161
rect 954 2158 1198 2161
rect 1266 2158 1278 2161
rect 1330 2158 1358 2161
rect 1362 2158 1406 2161
rect 1450 2158 1654 2161
rect 1658 2158 1702 2161
rect 1770 2158 1870 2161
rect 1922 2158 1966 2161
rect 1970 2158 2006 2161
rect 2098 2158 2102 2161
rect 2106 2158 2142 2161
rect 2146 2158 2174 2161
rect 2178 2158 2206 2161
rect 2250 2158 2254 2161
rect 2306 2158 2342 2161
rect 2370 2158 2374 2161
rect 2418 2158 2462 2161
rect 2474 2158 2598 2161
rect 2822 2161 2825 2168
rect 2934 2162 2937 2168
rect 2822 2158 2830 2161
rect 2914 2158 2926 2161
rect 2970 2158 3006 2161
rect 3070 2161 3073 2168
rect 3070 2158 3086 2161
rect 3154 2158 3230 2161
rect 3298 2158 3430 2161
rect 558 2152 561 2158
rect 18 2148 70 2151
rect 98 2148 118 2151
rect 170 2148 206 2151
rect 234 2148 249 2151
rect 338 2148 382 2151
rect 450 2148 510 2151
rect 602 2148 606 2151
rect 626 2148 726 2151
rect 754 2148 774 2151
rect 842 2148 902 2151
rect 1018 2148 1110 2151
rect 1114 2148 1118 2151
rect 1146 2148 1150 2151
rect 1194 2148 1222 2151
rect 1258 2148 1278 2151
rect 1298 2148 1334 2151
rect 1402 2148 1614 2151
rect 1618 2148 1630 2151
rect 1650 2148 1854 2151
rect 1858 2148 1990 2151
rect 1994 2148 2094 2151
rect 2098 2148 2246 2151
rect 2250 2148 2326 2151
rect 2330 2148 2606 2151
rect 2610 2148 2654 2151
rect 2690 2148 2750 2151
rect 2774 2151 2777 2158
rect 2754 2148 2777 2151
rect 2786 2148 2830 2151
rect 2834 2148 2862 2151
rect 2942 2151 2945 2158
rect 2898 2148 2945 2151
rect 2958 2148 3137 2151
rect 3154 2148 3158 2151
rect 3194 2148 3198 2151
rect 3218 2148 3222 2151
rect 3234 2148 3286 2151
rect 3338 2148 3342 2151
rect 3346 2148 3374 2151
rect 3590 2151 3594 2152
rect 3450 2148 3594 2151
rect 246 2142 249 2148
rect 798 2142 801 2148
rect 998 2142 1001 2148
rect 2958 2142 2961 2148
rect 82 2138 150 2141
rect 154 2138 158 2141
rect 178 2138 182 2141
rect 370 2138 414 2141
rect 418 2138 558 2141
rect 562 2138 569 2141
rect 578 2138 686 2141
rect 690 2138 774 2141
rect 810 2138 822 2141
rect 866 2138 886 2141
rect 890 2138 934 2141
rect 938 2138 982 2141
rect 1002 2138 1062 2141
rect 1114 2138 1126 2141
rect 1162 2138 1574 2141
rect 1626 2138 1638 2141
rect 1642 2138 1646 2141
rect 1786 2138 1790 2141
rect 1818 2138 1822 2141
rect 1842 2138 1846 2141
rect 1866 2138 1918 2141
rect 1962 2138 1966 2141
rect 1986 2138 2126 2141
rect 2130 2138 2190 2141
rect 2194 2138 2278 2141
rect 2282 2138 2302 2141
rect 2306 2138 2390 2141
rect 2394 2138 2414 2141
rect 2498 2138 2502 2141
rect 2530 2138 2534 2141
rect 2634 2138 2646 2141
rect 2670 2138 2697 2141
rect 2706 2138 2726 2141
rect 2842 2138 2846 2141
rect 2858 2138 2902 2141
rect 2906 2138 2958 2141
rect 2998 2138 3070 2141
rect 3134 2141 3137 2148
rect 3134 2138 3270 2141
rect 3274 2138 3486 2141
rect 566 2132 569 2138
rect 2670 2132 2673 2138
rect 2694 2132 2697 2138
rect 2998 2132 3001 2138
rect 18 2128 22 2131
rect 98 2128 174 2131
rect 178 2128 190 2131
rect 202 2128 214 2131
rect 218 2128 254 2131
rect 266 2128 310 2131
rect 346 2128 406 2131
rect 634 2128 646 2131
rect 658 2128 702 2131
rect 706 2128 710 2131
rect 714 2128 726 2131
rect 730 2128 758 2131
rect 762 2128 806 2131
rect 986 2128 1094 2131
rect 1098 2128 1294 2131
rect 1306 2128 1326 2131
rect 1506 2128 1734 2131
rect 1786 2128 1790 2131
rect 1818 2128 1918 2131
rect 1922 2128 2230 2131
rect 2242 2128 2254 2131
rect 2258 2128 2366 2131
rect 2578 2128 2630 2131
rect 2698 2128 2790 2131
rect 2874 2128 2910 2131
rect 2922 2128 2934 2131
rect 2938 2128 2990 2131
rect 3138 2128 3166 2131
rect 3290 2128 3294 2131
rect 3346 2128 3350 2131
rect 3354 2128 3406 2131
rect 3410 2128 3454 2131
rect 162 2118 342 2121
rect 354 2118 478 2121
rect 482 2118 550 2121
rect 570 2118 606 2121
rect 650 2118 686 2121
rect 922 2118 1086 2121
rect 1106 2118 1110 2121
rect 1210 2118 1246 2121
rect 1258 2118 1318 2121
rect 1514 2118 1574 2121
rect 1586 2118 1662 2121
rect 1762 2118 1870 2121
rect 1898 2118 1974 2121
rect 2018 2118 2070 2121
rect 2074 2118 2110 2121
rect 2114 2118 2326 2121
rect 2330 2118 2422 2121
rect 2426 2118 2462 2121
rect 2586 2118 2830 2121
rect 2866 2118 3030 2121
rect 3034 2118 3073 2121
rect 3082 2118 3262 2121
rect 3266 2118 3382 2121
rect 130 2108 326 2111
rect 458 2108 462 2111
rect 466 2108 518 2111
rect 522 2108 574 2111
rect 762 2108 870 2111
rect 1074 2108 1278 2111
rect 1282 2108 1286 2111
rect 1306 2108 1606 2111
rect 1614 2108 1750 2111
rect 1866 2108 1958 2111
rect 2050 2108 2062 2111
rect 2186 2108 2214 2111
rect 2226 2108 2270 2111
rect 2282 2108 2286 2111
rect 2330 2108 2358 2111
rect 2362 2108 2646 2111
rect 2650 2108 2742 2111
rect 2754 2108 2846 2111
rect 2850 2108 2910 2111
rect 3070 2111 3073 2118
rect 3070 2108 3238 2111
rect 3266 2108 3302 2111
rect 3330 2108 3446 2111
rect 630 2102 633 2108
rect 750 2102 753 2108
rect 992 2103 994 2107
rect 998 2103 1001 2107
rect 1006 2103 1008 2107
rect 242 2098 382 2101
rect 386 2098 454 2101
rect 594 2098 622 2101
rect 802 2098 838 2101
rect 1234 2098 1262 2101
rect 1338 2098 1438 2101
rect 1466 2098 1545 2101
rect 1614 2101 1617 2108
rect 2024 2103 2026 2107
rect 2030 2103 2033 2107
rect 2038 2103 2040 2107
rect 3040 2103 3042 2107
rect 3046 2103 3049 2107
rect 3054 2103 3056 2107
rect 1554 2098 1617 2101
rect 1650 2098 1726 2101
rect 1754 2098 1806 2101
rect 1818 2098 1846 2101
rect 1858 2098 1862 2101
rect 1890 2098 1926 2101
rect 2178 2098 2214 2101
rect 2234 2098 2342 2101
rect 2354 2098 2478 2101
rect 2514 2098 2534 2101
rect 2610 2098 2718 2101
rect 2722 2098 2742 2101
rect 2746 2098 2798 2101
rect 2834 2098 3030 2101
rect 3218 2098 3358 2101
rect 3362 2098 3390 2101
rect 3590 2101 3594 2102
rect 3490 2098 3594 2101
rect 910 2092 913 2098
rect 138 2088 166 2091
rect 186 2088 238 2091
rect 306 2088 470 2091
rect 522 2088 526 2091
rect 554 2088 758 2091
rect 770 2088 782 2091
rect 786 2088 790 2091
rect 826 2088 838 2091
rect 954 2088 1038 2091
rect 1050 2088 1070 2091
rect 1106 2088 1142 2091
rect 1202 2088 1206 2091
rect 1210 2088 1214 2091
rect 1226 2088 1286 2091
rect 1290 2088 1326 2091
rect 1330 2088 1334 2091
rect 1338 2088 1358 2091
rect 1362 2088 1366 2091
rect 1370 2088 1382 2091
rect 1386 2088 1390 2091
rect 1394 2088 1430 2091
rect 1434 2088 1454 2091
rect 1458 2088 1486 2091
rect 1542 2091 1545 2098
rect 1542 2088 1630 2091
rect 1722 2088 2606 2091
rect 2714 2088 2790 2091
rect 2794 2088 2894 2091
rect 2898 2088 2934 2091
rect 2938 2088 2966 2091
rect 3058 2088 3078 2091
rect 3114 2088 3182 2091
rect 266 2078 278 2081
rect 314 2078 318 2081
rect 346 2078 422 2081
rect 442 2078 625 2081
rect 634 2078 638 2081
rect 690 2078 694 2081
rect 754 2078 854 2081
rect 930 2078 934 2081
rect 1034 2078 1054 2081
rect 1066 2078 1118 2081
rect 1178 2078 1262 2081
rect 1394 2078 1398 2081
rect 1498 2078 1590 2081
rect 1686 2081 1689 2088
rect 1618 2078 1689 2081
rect 1770 2078 1822 2081
rect 1882 2078 1910 2081
rect 2066 2078 2150 2081
rect 2202 2078 2206 2081
rect 2226 2078 2238 2081
rect 2298 2078 2310 2081
rect 2346 2078 2382 2081
rect 2394 2078 2398 2081
rect 2410 2078 2414 2081
rect 2442 2078 2446 2081
rect 2490 2078 2502 2081
rect 2522 2078 2558 2081
rect 2738 2078 2758 2081
rect 2890 2078 2902 2081
rect 2946 2078 2974 2081
rect 3050 2078 3070 2081
rect 3090 2078 3102 2081
rect 3262 2081 3265 2088
rect 3262 2078 3366 2081
rect 86 2072 89 2078
rect 50 2068 70 2071
rect 166 2071 169 2078
rect 622 2072 625 2078
rect 1926 2072 1929 2078
rect 2166 2072 2169 2078
rect 90 2068 169 2071
rect 250 2068 262 2071
rect 274 2068 278 2071
rect 322 2068 526 2071
rect 530 2068 534 2071
rect 554 2068 606 2071
rect 626 2068 638 2071
rect 682 2068 710 2071
rect 802 2068 894 2071
rect 930 2068 998 2071
rect 1002 2068 1046 2071
rect 1050 2068 1262 2071
rect 1282 2068 1302 2071
rect 1314 2068 1318 2071
rect 1330 2068 1422 2071
rect 1570 2068 1710 2071
rect 1778 2068 1782 2071
rect 1946 2068 1998 2071
rect 2010 2068 2014 2071
rect 2058 2068 2094 2071
rect 2242 2068 2246 2071
rect 2290 2068 2294 2071
rect 2386 2068 2606 2071
rect 2678 2071 2681 2078
rect 2610 2068 2742 2071
rect 2782 2071 2785 2078
rect 3134 2072 3137 2078
rect 3150 2072 3153 2078
rect 3198 2072 3201 2078
rect 2778 2068 2785 2071
rect 2914 2068 2918 2071
rect 2922 2068 2929 2071
rect 3042 2068 3062 2071
rect 3074 2068 3094 2071
rect 3242 2068 3326 2071
rect 3354 2068 3374 2071
rect 3590 2071 3594 2072
rect 3562 2068 3594 2071
rect 74 2058 78 2061
rect 198 2061 201 2068
rect 146 2058 201 2061
rect 394 2058 494 2061
rect 498 2058 550 2061
rect 594 2058 614 2061
rect 658 2058 742 2061
rect 746 2058 838 2061
rect 866 2058 902 2061
rect 906 2058 982 2061
rect 1058 2058 1062 2061
rect 1098 2058 1606 2061
rect 1682 2058 1694 2061
rect 1726 2061 1729 2068
rect 1886 2062 1889 2068
rect 2318 2062 2321 2068
rect 1726 2058 1766 2061
rect 1850 2058 1878 2061
rect 1910 2058 2086 2061
rect 2098 2058 2102 2061
rect 2138 2058 2142 2061
rect 2170 2058 2174 2061
rect 2386 2058 2390 2061
rect 2402 2058 2486 2061
rect 2682 2058 2766 2061
rect 2786 2058 3318 2061
rect 3462 2061 3465 2068
rect 3370 2058 3433 2061
rect 3462 2058 3542 2061
rect 18 2048 22 2051
rect 66 2048 94 2051
rect 98 2048 758 2051
rect 778 2048 889 2051
rect 914 2048 918 2051
rect 946 2048 950 2051
rect 982 2051 985 2058
rect 1910 2052 1913 2058
rect 2190 2052 2193 2058
rect 2302 2052 2305 2058
rect 3430 2052 3433 2058
rect 982 2048 1110 2051
rect 1114 2048 1142 2051
rect 1146 2048 1166 2051
rect 1250 2048 1398 2051
rect 1570 2048 1574 2051
rect 1634 2048 1774 2051
rect 1858 2048 1862 2051
rect 1898 2048 1902 2051
rect 1946 2048 1998 2051
rect 2058 2048 2062 2051
rect 2130 2048 2134 2051
rect 2218 2048 2262 2051
rect 2346 2048 2350 2051
rect 2370 2048 2398 2051
rect 2434 2048 2462 2051
rect 2690 2048 2718 2051
rect 2762 2048 2814 2051
rect 2818 2048 2902 2051
rect 2922 2048 2977 2051
rect 2986 2048 3038 2051
rect 3058 2048 3078 2051
rect 3186 2048 3222 2051
rect 3354 2048 3358 2051
rect 3590 2051 3594 2052
rect 3562 2048 3594 2051
rect 886 2042 889 2048
rect 10 2038 46 2041
rect 50 2038 150 2041
rect 154 2038 262 2041
rect 354 2038 446 2041
rect 450 2038 598 2041
rect 602 2038 606 2041
rect 610 2038 654 2041
rect 666 2038 686 2041
rect 714 2038 718 2041
rect 834 2038 846 2041
rect 1014 2038 1030 2041
rect 1066 2038 1078 2041
rect 1202 2038 1254 2041
rect 1414 2041 1417 2048
rect 1502 2042 1505 2048
rect 1282 2038 1417 2041
rect 1442 2038 1502 2041
rect 1514 2038 1638 2041
rect 1642 2038 1694 2041
rect 1698 2038 1854 2041
rect 1858 2038 1982 2041
rect 1986 2038 2038 2041
rect 2042 2038 2070 2041
rect 2074 2038 2102 2041
rect 2118 2041 2121 2048
rect 2414 2042 2417 2048
rect 2486 2042 2489 2048
rect 2590 2042 2593 2048
rect 2654 2042 2657 2048
rect 2118 2038 2142 2041
rect 2162 2038 2198 2041
rect 2258 2038 2286 2041
rect 2314 2038 2406 2041
rect 2446 2038 2454 2041
rect 2458 2038 2478 2041
rect 2750 2041 2753 2048
rect 2722 2038 2753 2041
rect 2770 2038 2790 2041
rect 2810 2038 2942 2041
rect 2974 2041 2977 2048
rect 2974 2038 2998 2041
rect 3010 2038 3014 2041
rect 3210 2038 3294 2041
rect 1014 2032 1017 2038
rect 3126 2032 3129 2038
rect 82 2028 118 2031
rect 178 2028 302 2031
rect 466 2028 502 2031
rect 514 2028 694 2031
rect 746 2028 758 2031
rect 842 2028 1006 2031
rect 1026 2028 1078 2031
rect 1090 2028 1406 2031
rect 1418 2028 1598 2031
rect 1610 2028 1678 2031
rect 1682 2028 1734 2031
rect 1754 2028 1822 2031
rect 1842 2028 2478 2031
rect 2482 2028 2862 2031
rect 2874 2028 2878 2031
rect 2898 2028 2950 2031
rect 2954 2028 2966 2031
rect 250 2018 1646 2021
rect 1666 2018 1734 2021
rect 1778 2018 1782 2021
rect 1914 2018 1934 2021
rect 1946 2018 1950 2021
rect 1962 2018 1966 2021
rect 2106 2018 2294 2021
rect 2298 2018 2502 2021
rect 2506 2018 2534 2021
rect 2538 2018 2590 2021
rect 2602 2018 2654 2021
rect 2818 2018 2878 2021
rect 2922 2018 2942 2021
rect 2962 2018 3142 2021
rect 3402 2018 3494 2021
rect 3498 2018 3526 2021
rect 178 2008 262 2011
rect 426 2008 430 2011
rect 514 2008 526 2011
rect 618 2008 654 2011
rect 946 2008 1406 2011
rect 1602 2008 1678 2011
rect 1698 2008 1702 2011
rect 1874 2008 1918 2011
rect 1970 2008 2414 2011
rect 2442 2008 2446 2011
rect 2450 2008 2494 2011
rect 2514 2008 2518 2011
rect 2562 2008 2886 2011
rect 2890 2008 3054 2011
rect 3090 2008 3118 2011
rect 3122 2008 3238 2011
rect 3474 2008 3502 2011
rect 480 2003 482 2007
rect 486 2003 489 2007
rect 494 2003 496 2007
rect 1512 2003 1514 2007
rect 1518 2003 1521 2007
rect 1526 2003 1528 2007
rect 1934 2002 1937 2008
rect 1950 2002 1953 2008
rect 2536 2003 2538 2007
rect 2542 2003 2545 2007
rect 2550 2003 2552 2007
rect 218 1998 374 2001
rect 378 1998 462 2001
rect 506 1998 534 2001
rect 546 1998 1094 2001
rect 1266 1998 1310 2001
rect 1346 1998 1374 2001
rect 1442 1998 1478 2001
rect 1538 1998 1542 2001
rect 1546 1998 1606 2001
rect 1634 1998 1662 2001
rect 1714 1998 1782 2001
rect 1794 1998 1926 2001
rect 2146 1998 2422 2001
rect 2426 1998 2430 2001
rect 2450 1998 2518 2001
rect 2682 1998 2686 2001
rect 2898 1998 2990 2001
rect 3114 1998 3198 2001
rect 98 1988 230 1991
rect 290 1988 302 1991
rect 306 1988 358 1991
rect 378 1988 422 1991
rect 434 1988 470 1991
rect 478 1988 566 1991
rect 586 1988 590 1991
rect 626 1988 646 1991
rect 658 1988 662 1991
rect 674 1988 734 1991
rect 770 1988 774 1991
rect 794 1988 798 1991
rect 890 1988 950 1991
rect 962 1988 1046 1991
rect 1170 1988 1222 1991
rect 1274 1988 1286 1991
rect 1298 1988 2462 1991
rect 2466 1988 2734 1991
rect 2746 1988 2750 1991
rect 2762 1988 2838 1991
rect 2866 1988 2870 1991
rect 2914 1988 2926 1991
rect 2978 1988 3118 1991
rect 3138 1988 3230 1991
rect 3418 1988 3486 1991
rect 478 1982 481 1988
rect 266 1978 294 1981
rect 314 1978 318 1981
rect 418 1978 430 1981
rect 442 1978 478 1981
rect 530 1978 534 1981
rect 554 1978 694 1981
rect 730 1978 734 1981
rect 770 1978 910 1981
rect 962 1978 1022 1981
rect 1154 1978 1174 1981
rect 1194 1978 1270 1981
rect 1274 1978 1542 1981
rect 1682 1978 1726 1981
rect 1778 1978 1830 1981
rect 1850 1978 1878 1981
rect 2002 1978 2206 1981
rect 2258 1978 2462 1981
rect 2466 1978 2694 1981
rect 2698 1978 2878 1981
rect 2970 1978 3150 1981
rect 3154 1978 3174 1981
rect 166 1972 169 1978
rect 242 1968 558 1971
rect 570 1968 774 1971
rect 786 1968 798 1971
rect 930 1968 966 1971
rect 1022 1971 1025 1978
rect 1022 1968 1038 1971
rect 1102 1971 1105 1978
rect 1050 1968 1105 1971
rect 1122 1968 1126 1971
rect 1130 1968 1238 1971
rect 1250 1968 1462 1971
rect 1482 1968 1686 1971
rect 1746 1968 1750 1971
rect 1958 1971 1961 1978
rect 1958 1968 2046 1971
rect 2090 1968 2094 1971
rect 2162 1968 2206 1971
rect 2282 1968 2710 1971
rect 2714 1968 2950 1971
rect 3010 1968 3014 1971
rect 3034 1968 3070 1971
rect 3298 1968 3430 1971
rect 3474 1968 3486 1971
rect 3518 1971 3521 1978
rect 3590 1971 3594 1972
rect 3518 1968 3594 1971
rect 118 1962 121 1968
rect 1718 1962 1721 1968
rect 1726 1962 1729 1968
rect 1862 1962 1865 1968
rect 74 1958 94 1961
rect 162 1958 174 1961
rect 194 1958 438 1961
rect 466 1958 526 1961
rect 530 1958 582 1961
rect 586 1958 606 1961
rect 650 1958 662 1961
rect 682 1958 1030 1961
rect 1034 1958 1086 1961
rect 1090 1958 1326 1961
rect 1338 1958 1342 1961
rect 1466 1958 1470 1961
rect 1490 1958 1518 1961
rect 1546 1958 1590 1961
rect 1626 1958 1654 1961
rect 1666 1958 1694 1961
rect 1826 1958 1838 1961
rect 1930 1958 1934 1961
rect 2110 1961 2113 1968
rect 1954 1958 2113 1961
rect 2154 1958 2174 1961
rect 2234 1958 2262 1961
rect 2274 1958 2318 1961
rect 2366 1958 2374 1961
rect 2378 1958 2390 1961
rect 2682 1958 2686 1961
rect 2730 1958 2918 1961
rect 2930 1958 2958 1961
rect 3126 1961 3129 1968
rect 2966 1958 3129 1961
rect 3162 1958 3190 1961
rect 3246 1961 3249 1968
rect 3202 1958 3249 1961
rect 3266 1958 3270 1961
rect 3282 1958 3302 1961
rect 3306 1958 3334 1961
rect 3338 1958 3342 1961
rect 3418 1958 3502 1961
rect 638 1952 641 1958
rect 1358 1952 1361 1958
rect 42 1948 86 1951
rect 130 1948 134 1951
rect 154 1948 206 1951
rect 218 1948 278 1951
rect 290 1948 334 1951
rect 338 1948 382 1951
rect 402 1948 430 1951
rect 450 1948 582 1951
rect 586 1948 606 1951
rect 610 1948 614 1951
rect 650 1948 710 1951
rect 714 1948 758 1951
rect 762 1948 854 1951
rect 906 1948 918 1951
rect 946 1948 966 1951
rect 1018 1948 1070 1951
rect 1138 1948 1166 1951
rect 1178 1948 1182 1951
rect 1298 1948 1302 1951
rect 1330 1948 1342 1951
rect 1386 1948 1406 1951
rect 1410 1948 1414 1951
rect 1442 1948 1558 1951
rect 1666 1948 1670 1951
rect 1710 1948 1774 1951
rect 1786 1948 1838 1951
rect 1850 1948 1854 1951
rect 1866 1948 1942 1951
rect 1946 1948 1998 1951
rect 2002 1948 2006 1951
rect 2034 1948 2078 1951
rect 2122 1948 2358 1951
rect 2386 1948 2390 1951
rect 2486 1951 2489 1958
rect 2482 1948 2489 1951
rect 2606 1952 2609 1958
rect 2658 1948 2766 1951
rect 2778 1948 2798 1951
rect 2802 1948 2822 1951
rect 2850 1948 2918 1951
rect 2966 1951 2969 1958
rect 2930 1948 2969 1951
rect 3142 1951 3145 1958
rect 3010 1948 3105 1951
rect 3142 1948 3190 1951
rect 3194 1948 3206 1951
rect 3266 1948 3270 1951
rect 3358 1951 3361 1958
rect 3282 1948 3361 1951
rect 3390 1951 3393 1958
rect 3390 1948 3446 1951
rect 3482 1948 3518 1951
rect 3590 1951 3594 1952
rect 3562 1948 3594 1951
rect 174 1942 177 1948
rect 10 1938 30 1941
rect 34 1938 94 1941
rect 98 1938 118 1941
rect 282 1938 350 1941
rect 354 1938 390 1941
rect 478 1938 526 1941
rect 562 1938 630 1941
rect 634 1938 646 1941
rect 666 1938 766 1941
rect 778 1938 822 1941
rect 914 1938 942 1941
rect 978 1938 982 1941
rect 1106 1938 1142 1941
rect 1146 1938 1190 1941
rect 1250 1938 1254 1941
rect 1422 1941 1425 1948
rect 1290 1938 1425 1941
rect 1434 1938 1446 1941
rect 1498 1938 1542 1941
rect 1554 1938 1558 1941
rect 1578 1938 1582 1941
rect 1626 1938 1641 1941
rect 1650 1938 1686 1941
rect 1710 1941 1713 1948
rect 2094 1942 2097 1948
rect 3102 1942 3105 1948
rect 1690 1938 1713 1941
rect 1722 1938 1742 1941
rect 1762 1938 1966 1941
rect 2138 1938 2166 1941
rect 2170 1938 2230 1941
rect 2238 1938 2310 1941
rect 2322 1938 2334 1941
rect 2530 1938 2550 1941
rect 2642 1938 2702 1941
rect 2706 1938 2766 1941
rect 2858 1938 2870 1941
rect 2914 1938 2918 1941
rect 2938 1938 2942 1941
rect 2962 1938 2985 1941
rect 3050 1938 3054 1941
rect 3202 1938 3206 1941
rect 3234 1938 3302 1941
rect 3458 1938 3518 1941
rect 478 1932 481 1938
rect 766 1932 769 1938
rect 1566 1932 1569 1938
rect 1638 1932 1641 1938
rect 1974 1932 1977 1938
rect 2238 1932 2241 1938
rect 2982 1932 2985 1938
rect 158 1928 166 1931
rect 170 1928 230 1931
rect 530 1928 534 1931
rect 538 1928 542 1931
rect 650 1928 678 1931
rect 698 1928 742 1931
rect 746 1928 750 1931
rect 890 1928 942 1931
rect 978 1928 1206 1931
rect 1298 1928 1302 1931
rect 1314 1928 1366 1931
rect 1386 1928 1390 1931
rect 1466 1928 1534 1931
rect 1546 1928 1550 1931
rect 1578 1928 1590 1931
rect 1602 1928 1630 1931
rect 1642 1928 1742 1931
rect 1770 1928 1774 1931
rect 1802 1928 1806 1931
rect 1826 1928 1870 1931
rect 1890 1928 1894 1931
rect 1906 1928 1918 1931
rect 1930 1928 1942 1931
rect 2042 1928 2054 1931
rect 2090 1928 2150 1931
rect 2154 1928 2182 1931
rect 2186 1928 2214 1931
rect 2258 1928 2270 1931
rect 2298 1928 2326 1931
rect 2482 1928 2566 1931
rect 2662 1928 2814 1931
rect 2882 1928 2950 1931
rect 3070 1931 3073 1938
rect 3070 1928 3158 1931
rect 3162 1928 3222 1931
rect 3242 1928 3270 1931
rect 3322 1928 3382 1931
rect 106 1918 254 1921
rect 290 1918 406 1921
rect 474 1918 638 1921
rect 646 1918 1758 1921
rect 1770 1918 1774 1921
rect 1782 1921 1785 1928
rect 1782 1918 1814 1921
rect 1866 1918 1870 1921
rect 1878 1921 1881 1928
rect 2374 1922 2377 1928
rect 2662 1922 2665 1928
rect 1878 1918 1910 1921
rect 1946 1918 1982 1921
rect 1986 1918 2030 1921
rect 2042 1918 2094 1921
rect 2106 1918 2238 1921
rect 2242 1918 2353 1921
rect 2738 1918 2742 1921
rect 2754 1918 2774 1921
rect 2778 1918 2785 1921
rect 2794 1918 3278 1921
rect 122 1908 214 1911
rect 226 1908 310 1911
rect 314 1908 502 1911
rect 530 1908 574 1911
rect 646 1911 649 1918
rect 1838 1912 1841 1918
rect 1846 1912 1849 1918
rect 634 1908 649 1911
rect 746 1908 774 1911
rect 866 1908 878 1911
rect 1058 1908 1214 1911
rect 1226 1908 1286 1911
rect 1362 1908 1430 1911
rect 1506 1908 1665 1911
rect 1714 1908 1782 1911
rect 1802 1908 1822 1911
rect 1858 1908 1990 1911
rect 2050 1908 2062 1911
rect 2082 1908 2118 1911
rect 2154 1908 2158 1911
rect 2170 1908 2190 1911
rect 2210 1908 2246 1911
rect 2350 1911 2353 1918
rect 2350 1908 2454 1911
rect 2458 1908 2486 1911
rect 2498 1908 2574 1911
rect 2610 1908 2710 1911
rect 2762 1908 2854 1911
rect 2914 1908 2918 1911
rect 2970 1908 3014 1911
rect 3122 1908 3214 1911
rect 694 1902 697 1908
rect 992 1903 994 1907
rect 998 1903 1001 1907
rect 1006 1903 1008 1907
rect 1662 1902 1665 1908
rect 2024 1903 2026 1907
rect 2030 1903 2033 1907
rect 2038 1903 2040 1907
rect 3040 1903 3042 1907
rect 3046 1903 3049 1907
rect 3054 1903 3056 1907
rect 98 1898 142 1901
rect 202 1898 318 1901
rect 338 1898 382 1901
rect 386 1898 414 1901
rect 426 1898 430 1901
rect 458 1898 638 1901
rect 682 1898 686 1901
rect 746 1898 870 1901
rect 930 1898 934 1901
rect 938 1898 974 1901
rect 1014 1898 1614 1901
rect 1666 1898 1678 1901
rect 1706 1898 1798 1901
rect 1810 1898 1822 1901
rect 1834 1898 1993 1901
rect 2138 1898 2158 1901
rect 2202 1898 2214 1901
rect 2226 1898 2494 1901
rect 2618 1898 2622 1901
rect 2626 1898 2974 1901
rect 2994 1898 3022 1901
rect 3066 1898 3230 1901
rect 3234 1898 3502 1901
rect 3514 1898 3526 1901
rect 1014 1891 1017 1898
rect 1990 1892 1993 1898
rect 146 1888 1017 1891
rect 1114 1888 1230 1891
rect 1290 1888 1318 1891
rect 1394 1888 1494 1891
rect 1554 1888 1862 1891
rect 1866 1888 1937 1891
rect 102 1881 105 1888
rect 1934 1882 1937 1888
rect 2010 1888 2038 1891
rect 2050 1888 2214 1891
rect 2234 1888 2238 1891
rect 2250 1888 2254 1891
rect 2298 1888 2302 1891
rect 2322 1888 2326 1891
rect 2410 1888 2486 1891
rect 2698 1888 2718 1891
rect 2842 1888 2857 1891
rect 2874 1888 2894 1891
rect 2930 1888 3078 1891
rect 3118 1888 3126 1891
rect 3146 1888 3230 1891
rect 3330 1888 3374 1891
rect 3378 1888 3478 1891
rect 18 1878 105 1881
rect 210 1878 222 1881
rect 490 1878 510 1881
rect 562 1878 590 1881
rect 618 1878 630 1881
rect 642 1878 798 1881
rect 826 1878 982 1881
rect 1002 1878 1054 1881
rect 1058 1878 1086 1881
rect 1098 1878 1150 1881
rect 1162 1878 1166 1881
rect 1186 1878 1225 1881
rect 1234 1878 1278 1881
rect 1434 1878 1502 1881
rect 1658 1878 1926 1881
rect 1990 1881 1993 1888
rect 1990 1878 2022 1881
rect 2210 1878 2334 1881
rect 2354 1878 2590 1881
rect 2654 1881 2657 1888
rect 2634 1878 2657 1881
rect 2674 1878 2678 1881
rect 2698 1878 2710 1881
rect 2842 1878 2846 1881
rect 2854 1881 2857 1888
rect 3118 1882 3121 1888
rect 2854 1878 2918 1881
rect 3226 1878 3318 1881
rect 3514 1878 3526 1881
rect 34 1868 46 1871
rect 90 1868 110 1871
rect 210 1868 222 1871
rect 274 1868 366 1871
rect 722 1868 750 1871
rect 754 1868 766 1871
rect 770 1868 830 1871
rect 834 1868 862 1871
rect 866 1868 886 1871
rect 922 1868 934 1871
rect 994 1868 998 1871
rect 1090 1868 1174 1871
rect 1210 1868 1214 1871
rect 1222 1871 1225 1878
rect 1318 1872 1321 1878
rect 1222 1868 1254 1871
rect 1258 1868 1278 1871
rect 1370 1868 1374 1871
rect 1442 1868 1446 1871
rect 1458 1868 1486 1871
rect 1490 1868 1582 1871
rect 1638 1871 1641 1878
rect 2686 1872 2689 1878
rect 1594 1868 1641 1871
rect 1650 1868 1662 1871
rect 1674 1868 1886 1871
rect 1922 1868 2006 1871
rect 2010 1868 2129 1871
rect 2146 1868 2174 1871
rect 2242 1868 2342 1871
rect 2386 1868 2454 1871
rect 2458 1868 2622 1871
rect 2626 1868 2630 1871
rect 2658 1868 2670 1871
rect 2706 1868 2710 1871
rect 2778 1868 2830 1871
rect 2834 1868 2870 1871
rect 2906 1868 2926 1871
rect 2930 1868 2966 1871
rect 3002 1868 3006 1871
rect 3082 1868 3086 1871
rect 3154 1868 3254 1871
rect 3402 1868 3454 1871
rect 3590 1871 3594 1872
rect 3546 1868 3594 1871
rect 582 1862 585 1868
rect 614 1862 617 1868
rect 34 1858 230 1861
rect 306 1858 318 1861
rect 322 1858 334 1861
rect 626 1858 646 1861
rect 770 1858 774 1861
rect 818 1858 838 1861
rect 930 1858 1374 1861
rect 1402 1858 1422 1861
rect 1450 1858 1486 1861
rect 1498 1858 1518 1861
rect 1538 1858 1598 1861
rect 1614 1858 1622 1861
rect 1642 1858 1670 1861
rect 1690 1858 1694 1861
rect 1706 1858 1710 1861
rect 1730 1858 1734 1861
rect 1754 1858 1758 1861
rect 1818 1858 1870 1861
rect 1930 1858 2118 1861
rect 2126 1861 2129 1868
rect 3222 1862 3225 1868
rect 2126 1858 2142 1861
rect 2162 1858 2270 1861
rect 2282 1858 2286 1861
rect 2298 1858 2366 1861
rect 2530 1858 2593 1861
rect 2666 1858 2734 1861
rect 2842 1858 2846 1861
rect 2946 1858 2990 1861
rect 3010 1858 3014 1861
rect 3082 1858 3102 1861
rect 3130 1858 3206 1861
rect 3234 1858 3262 1861
rect 3410 1859 3454 1861
rect 3410 1858 3457 1859
rect 30 1852 33 1858
rect 98 1848 102 1851
rect 170 1848 174 1851
rect 246 1851 249 1858
rect 246 1848 446 1851
rect 466 1848 518 1851
rect 530 1848 534 1851
rect 538 1848 590 1851
rect 698 1848 734 1851
rect 758 1851 761 1858
rect 758 1848 774 1851
rect 814 1851 817 1858
rect 1614 1852 1617 1858
rect 1886 1852 1889 1858
rect 794 1848 817 1851
rect 962 1848 966 1851
rect 1034 1848 1057 1851
rect 1130 1848 1262 1851
rect 1354 1848 1454 1851
rect 1466 1848 1542 1851
rect 1594 1848 1598 1851
rect 1626 1848 1670 1851
rect 1714 1848 1718 1851
rect 1770 1848 1806 1851
rect 1810 1848 1814 1851
rect 1834 1848 1862 1851
rect 1874 1848 1878 1851
rect 1914 1848 1974 1851
rect 1986 1848 1990 1851
rect 2002 1848 2006 1851
rect 2018 1848 2022 1851
rect 2082 1848 2270 1851
rect 2278 1848 2286 1851
rect 2290 1848 2302 1851
rect 2330 1848 2334 1851
rect 2490 1848 2582 1851
rect 2590 1851 2593 1858
rect 2998 1852 3001 1858
rect 3118 1852 3121 1858
rect 2590 1848 2622 1851
rect 2746 1848 2758 1851
rect 2826 1848 2958 1851
rect 3042 1848 3118 1851
rect 3154 1848 3158 1851
rect 3206 1851 3209 1858
rect 3206 1848 3254 1851
rect 3258 1848 3286 1851
rect 3402 1848 3406 1851
rect 3590 1851 3594 1852
rect 3562 1848 3594 1851
rect 590 1842 593 1848
rect 82 1838 150 1841
rect 298 1838 350 1841
rect 354 1838 374 1841
rect 378 1838 398 1841
rect 1054 1841 1057 1848
rect 1342 1842 1345 1848
rect 1054 1838 1134 1841
rect 1146 1838 1214 1841
rect 1226 1838 1294 1841
rect 1394 1838 1398 1841
rect 1506 1838 1598 1841
rect 1894 1841 1897 1848
rect 1610 1838 1897 1841
rect 1906 1838 2070 1841
rect 2098 1838 2345 1841
rect 2434 1838 2998 1841
rect 3002 1838 3174 1841
rect 3178 1838 3542 1841
rect 130 1828 222 1831
rect 518 1831 521 1838
rect 2342 1832 2345 1838
rect 362 1828 521 1831
rect 530 1828 550 1831
rect 594 1828 926 1831
rect 938 1828 1214 1831
rect 1250 1828 1334 1831
rect 1338 1828 1438 1831
rect 1442 1828 1617 1831
rect 1634 1828 1638 1831
rect 1674 1828 1814 1831
rect 1866 1828 1894 1831
rect 1914 1828 1918 1831
rect 1938 1828 1990 1831
rect 1994 1828 2262 1831
rect 2274 1828 2334 1831
rect 2346 1828 2558 1831
rect 2602 1828 2614 1831
rect 2650 1828 2702 1831
rect 2714 1828 2750 1831
rect 2794 1828 2814 1831
rect 2818 1828 2854 1831
rect 2858 1828 3510 1831
rect 3590 1831 3594 1832
rect 3514 1828 3594 1831
rect 310 1822 313 1828
rect 426 1818 438 1821
rect 442 1818 606 1821
rect 914 1818 950 1821
rect 978 1818 1222 1821
rect 1298 1818 1422 1821
rect 1426 1818 1454 1821
rect 1530 1818 1542 1821
rect 1570 1818 1606 1821
rect 1614 1821 1617 1828
rect 1614 1818 2430 1821
rect 2442 1818 2446 1821
rect 2450 1818 2558 1821
rect 2586 1818 2670 1821
rect 2722 1818 2902 1821
rect 2938 1818 3102 1821
rect 3146 1818 3150 1821
rect 3250 1818 3278 1821
rect 3330 1818 3438 1821
rect 66 1808 326 1811
rect 650 1808 806 1811
rect 810 1808 958 1811
rect 1098 1808 1225 1811
rect 1282 1808 1366 1811
rect 1402 1808 1414 1811
rect 1426 1808 1446 1811
rect 1466 1808 1470 1811
rect 1546 1808 1598 1811
rect 1610 1808 1646 1811
rect 1690 1808 1766 1811
rect 1786 1808 1790 1811
rect 1818 1808 1862 1811
rect 1874 1808 1926 1811
rect 1938 1808 2310 1811
rect 2338 1808 2401 1811
rect 2418 1808 2422 1811
rect 2562 1808 2630 1811
rect 2642 1808 2678 1811
rect 2770 1808 2934 1811
rect 3098 1808 3502 1811
rect 3590 1808 3594 1812
rect 480 1803 482 1807
rect 486 1803 489 1807
rect 494 1803 496 1807
rect 1222 1802 1225 1808
rect 1512 1803 1514 1807
rect 1518 1803 1521 1807
rect 1526 1803 1528 1807
rect 74 1798 294 1801
rect 410 1798 470 1801
rect 506 1798 598 1801
rect 762 1798 798 1801
rect 834 1798 926 1801
rect 1082 1798 1134 1801
rect 1138 1798 1174 1801
rect 1186 1798 1190 1801
rect 1226 1798 1270 1801
rect 1298 1798 1326 1801
rect 1338 1798 1470 1801
rect 1578 1798 1670 1801
rect 1682 1798 1742 1801
rect 1746 1798 1798 1801
rect 1802 1798 1958 1801
rect 1978 1798 1990 1801
rect 2074 1798 2078 1801
rect 2090 1798 2110 1801
rect 2398 1801 2401 1808
rect 2494 1802 2497 1808
rect 2536 1803 2538 1807
rect 2542 1803 2545 1807
rect 2550 1803 2552 1807
rect 2154 1798 2393 1801
rect 2398 1798 2414 1801
rect 2418 1798 2454 1801
rect 2586 1798 2598 1801
rect 2682 1798 2758 1801
rect 2770 1798 2790 1801
rect 2882 1798 3494 1801
rect 3590 1801 3593 1808
rect 3498 1798 3593 1801
rect 394 1788 566 1791
rect 778 1788 798 1791
rect 818 1788 958 1791
rect 1018 1788 1118 1791
rect 1194 1788 1654 1791
rect 1658 1788 2150 1791
rect 2194 1788 2198 1791
rect 2258 1788 2262 1791
rect 2274 1788 2278 1791
rect 2390 1791 2393 1798
rect 2654 1792 2657 1798
rect 2390 1788 2510 1791
rect 2514 1788 2606 1791
rect 2682 1788 2798 1791
rect 2802 1788 2934 1791
rect 3298 1788 3302 1791
rect 3366 1788 3390 1791
rect 3394 1788 3478 1791
rect 3590 1788 3594 1792
rect 254 1782 257 1788
rect 114 1778 142 1781
rect 530 1778 622 1781
rect 718 1778 905 1781
rect 914 1778 918 1781
rect 970 1778 1054 1781
rect 1090 1778 1126 1781
rect 1134 1781 1137 1788
rect 1134 1778 1254 1781
rect 1386 1778 1494 1781
rect 1506 1778 1510 1781
rect 1562 1778 1710 1781
rect 1722 1778 1734 1781
rect 1746 1778 1830 1781
rect 1930 1778 1934 1781
rect 1962 1778 1998 1781
rect 2002 1778 2222 1781
rect 2334 1781 2337 1788
rect 2226 1778 2366 1781
rect 2370 1778 2390 1781
rect 2570 1778 2670 1781
rect 2722 1778 2790 1781
rect 3230 1781 3233 1788
rect 3366 1782 3369 1788
rect 2946 1778 3233 1781
rect 3290 1778 3358 1781
rect 3410 1778 3430 1781
rect 3590 1781 3593 1788
rect 3562 1778 3593 1781
rect 718 1772 721 1778
rect 74 1768 166 1771
rect 210 1768 254 1771
rect 258 1768 262 1771
rect 362 1768 382 1771
rect 418 1768 438 1771
rect 458 1768 542 1771
rect 690 1768 702 1771
rect 706 1768 710 1771
rect 778 1768 822 1771
rect 902 1771 905 1778
rect 902 1768 918 1771
rect 922 1768 982 1771
rect 994 1768 1030 1771
rect 1062 1771 1065 1778
rect 1062 1768 1094 1771
rect 1138 1768 1326 1771
rect 1338 1768 1350 1771
rect 1362 1768 1534 1771
rect 1574 1768 1654 1771
rect 1714 1768 1774 1771
rect 1778 1768 1830 1771
rect 1842 1768 1870 1771
rect 1882 1768 1918 1771
rect 1922 1768 1950 1771
rect 1970 1768 2006 1771
rect 2010 1768 2094 1771
rect 2122 1768 2502 1771
rect 2506 1768 2654 1771
rect 2730 1768 2790 1771
rect 2794 1768 2830 1771
rect 2922 1768 3422 1771
rect 3590 1768 3594 1772
rect 62 1761 65 1768
rect 34 1758 86 1761
rect 110 1758 134 1761
rect 194 1758 270 1761
rect 274 1758 294 1761
rect 378 1758 662 1761
rect 666 1758 710 1761
rect 730 1758 1014 1761
rect 1042 1758 1046 1761
rect 1082 1758 1150 1761
rect 1154 1758 1158 1761
rect 1258 1758 1286 1761
rect 1346 1758 1350 1761
rect 1370 1758 1390 1761
rect 1442 1758 1446 1761
rect 1574 1761 1577 1768
rect 1498 1758 1577 1761
rect 1586 1758 1590 1761
rect 1626 1758 1638 1761
rect 1650 1758 1750 1761
rect 1778 1758 1854 1761
rect 1866 1758 1942 1761
rect 1962 1758 2054 1761
rect 2066 1758 2102 1761
rect 2114 1758 2118 1761
rect 2122 1758 2206 1761
rect 2210 1758 2230 1761
rect 2290 1758 2430 1761
rect 2458 1758 2694 1761
rect 2750 1758 2830 1761
rect 2834 1758 3006 1761
rect 3034 1758 3086 1761
rect 3114 1758 3182 1761
rect 3186 1758 3262 1761
rect 3590 1761 3593 1768
rect 3306 1758 3593 1761
rect 110 1752 113 1758
rect 158 1752 161 1758
rect 350 1752 353 1758
rect 2662 1752 2665 1758
rect 2750 1752 2753 1758
rect 42 1748 86 1751
rect 402 1748 422 1751
rect 466 1748 526 1751
rect 626 1748 662 1751
rect 674 1748 678 1751
rect 690 1748 702 1751
rect 722 1748 734 1751
rect 754 1748 774 1751
rect 906 1748 1022 1751
rect 1026 1748 1206 1751
rect 1266 1748 1270 1751
rect 1290 1748 1297 1751
rect 1306 1748 1310 1751
rect 1402 1748 1406 1751
rect 1418 1748 1422 1751
rect 1482 1748 1489 1751
rect 1522 1748 1542 1751
rect 1634 1748 1830 1751
rect 1842 1748 1846 1751
rect 1922 1748 1990 1751
rect 2042 1748 2118 1751
rect 2146 1748 2150 1751
rect 2202 1748 2214 1751
rect 2218 1748 2222 1751
rect 2258 1748 2278 1751
rect 2322 1748 2390 1751
rect 2410 1748 2438 1751
rect 2458 1748 2462 1751
rect 2518 1748 2526 1751
rect 2530 1748 2534 1751
rect 2578 1748 2598 1751
rect 2706 1748 2718 1751
rect 2722 1748 2750 1751
rect 2818 1748 2894 1751
rect 2898 1748 2966 1751
rect 2970 1748 2982 1751
rect 3066 1748 3070 1751
rect 3202 1748 3206 1751
rect 3210 1748 3254 1751
rect 3362 1748 3374 1751
rect 3378 1748 3438 1751
rect 3442 1748 3534 1751
rect 3590 1751 3594 1752
rect 3562 1748 3594 1751
rect 238 1742 241 1748
rect 26 1738 62 1741
rect 66 1738 78 1741
rect 122 1738 158 1741
rect 178 1738 198 1741
rect 282 1738 366 1741
rect 422 1738 430 1741
rect 434 1738 454 1741
rect 490 1738 494 1741
rect 538 1738 542 1741
rect 586 1738 606 1741
rect 610 1738 614 1741
rect 642 1738 646 1741
rect 658 1738 694 1741
rect 722 1738 766 1741
rect 778 1738 870 1741
rect 890 1738 945 1741
rect 970 1738 1030 1741
rect 1034 1738 1086 1741
rect 1114 1738 1134 1741
rect 1186 1738 1230 1741
rect 1250 1738 1278 1741
rect 1294 1741 1297 1748
rect 1366 1742 1369 1748
rect 1382 1742 1385 1748
rect 1486 1742 1489 1748
rect 1294 1738 1326 1741
rect 1402 1738 1422 1741
rect 1578 1738 1582 1741
rect 1590 1741 1593 1748
rect 1862 1742 1865 1748
rect 1590 1738 1606 1741
rect 1642 1738 1710 1741
rect 1730 1738 1734 1741
rect 1754 1738 1822 1741
rect 1834 1738 1838 1741
rect 1910 1741 1913 1748
rect 2254 1742 2257 1748
rect 2806 1742 2809 1748
rect 1910 1738 1926 1741
rect 2050 1738 2054 1741
rect 2106 1738 2126 1741
rect 2138 1738 2142 1741
rect 2162 1738 2182 1741
rect 2186 1738 2254 1741
rect 2274 1738 2302 1741
rect 2306 1738 2438 1741
rect 2594 1738 2670 1741
rect 2674 1738 2694 1741
rect 2698 1738 2726 1741
rect 2890 1738 2942 1741
rect 3074 1738 3086 1741
rect 3090 1738 3150 1741
rect 3234 1738 3238 1741
rect 3242 1738 3262 1741
rect 3266 1738 3294 1741
rect 3354 1738 3406 1741
rect 3418 1738 3422 1741
rect 3426 1738 3494 1741
rect 3530 1738 3534 1741
rect 230 1732 233 1738
rect 510 1732 513 1738
rect 942 1732 945 1738
rect 1110 1732 1113 1738
rect 10 1728 38 1731
rect 50 1728 174 1731
rect 242 1728 321 1731
rect 318 1722 321 1728
rect 410 1728 502 1731
rect 514 1728 790 1731
rect 794 1728 846 1731
rect 850 1728 918 1731
rect 930 1728 934 1731
rect 962 1728 1033 1731
rect 1042 1728 1054 1731
rect 1058 1728 1065 1731
rect 1130 1728 1201 1731
rect 1210 1728 1214 1731
rect 1274 1728 1278 1731
rect 1394 1728 1422 1731
rect 1426 1728 1526 1731
rect 1554 1728 1558 1731
rect 1578 1728 1590 1731
rect 1594 1728 1598 1731
rect 1610 1728 1638 1731
rect 1650 1728 1678 1731
rect 1706 1728 1710 1731
rect 1718 1728 1750 1731
rect 1786 1728 1798 1731
rect 1810 1728 1830 1731
rect 1850 1728 1886 1731
rect 1898 1728 1934 1731
rect 1994 1728 2022 1731
rect 2034 1728 2078 1731
rect 2114 1728 2126 1731
rect 2130 1728 2134 1731
rect 2170 1728 2286 1731
rect 2302 1728 2310 1731
rect 2314 1728 2358 1731
rect 2378 1728 2422 1731
rect 2578 1728 2646 1731
rect 2650 1728 2814 1731
rect 2838 1731 2841 1738
rect 2818 1728 2998 1731
rect 3002 1728 3110 1731
rect 3138 1728 3150 1731
rect 3154 1728 3206 1731
rect 3290 1728 3414 1731
rect 3418 1728 3473 1731
rect 3506 1728 3510 1731
rect 3590 1731 3594 1732
rect 3562 1728 3594 1731
rect 334 1722 337 1728
rect 106 1718 134 1721
rect 154 1718 310 1721
rect 442 1718 534 1721
rect 698 1718 702 1721
rect 882 1718 958 1721
rect 1030 1721 1033 1728
rect 962 1718 1025 1721
rect 1030 1718 1158 1721
rect 1162 1718 1190 1721
rect 1198 1721 1201 1728
rect 1318 1722 1321 1728
rect 1198 1718 1302 1721
rect 1362 1718 1454 1721
rect 1490 1718 1566 1721
rect 1650 1718 1654 1721
rect 1718 1721 1721 1728
rect 1674 1718 1721 1721
rect 1746 1718 1750 1721
rect 1770 1718 1774 1721
rect 1802 1718 1814 1721
rect 1826 1718 1846 1721
rect 1850 1718 1862 1721
rect 1874 1718 1918 1721
rect 1930 1718 2174 1721
rect 2202 1718 2278 1721
rect 2430 1721 2433 1728
rect 3470 1722 3473 1728
rect 2286 1718 2510 1721
rect 2514 1718 2574 1721
rect 2626 1718 2910 1721
rect 2946 1718 2950 1721
rect 2978 1718 3302 1721
rect 3482 1718 3518 1721
rect 3554 1718 3558 1721
rect 558 1712 561 1718
rect 590 1712 593 1718
rect 646 1712 649 1718
rect 34 1708 190 1711
rect 226 1708 238 1711
rect 378 1708 382 1711
rect 578 1708 582 1711
rect 658 1708 678 1711
rect 730 1708 742 1711
rect 818 1708 854 1711
rect 890 1708 910 1711
rect 930 1708 966 1711
rect 1022 1711 1025 1718
rect 1022 1708 1086 1711
rect 1098 1708 1102 1711
rect 1122 1708 1126 1711
rect 1138 1708 1166 1711
rect 1202 1708 1406 1711
rect 1442 1708 1502 1711
rect 1554 1708 1742 1711
rect 1754 1708 1870 1711
rect 1882 1708 1958 1711
rect 1986 1708 1998 1711
rect 2082 1708 2118 1711
rect 2130 1708 2166 1711
rect 2286 1711 2289 1718
rect 2178 1708 2289 1711
rect 2330 1708 2342 1711
rect 2354 1708 2390 1711
rect 2466 1708 2502 1711
rect 2562 1708 2678 1711
rect 2690 1708 2710 1711
rect 2778 1708 3030 1711
rect 3082 1708 3142 1711
rect 3146 1708 3198 1711
rect 3218 1708 3486 1711
rect 3530 1708 3542 1711
rect 992 1703 994 1707
rect 998 1703 1001 1707
rect 1006 1703 1008 1707
rect 2024 1703 2026 1707
rect 2030 1703 2033 1707
rect 2038 1703 2040 1707
rect 3040 1703 3042 1707
rect 3046 1703 3049 1707
rect 3054 1703 3056 1707
rect 82 1698 286 1701
rect 290 1698 478 1701
rect 538 1698 654 1701
rect 858 1698 910 1701
rect 914 1698 985 1701
rect 1034 1698 1158 1701
rect 1162 1698 1230 1701
rect 1330 1698 1478 1701
rect 1522 1698 1550 1701
rect 1634 1698 1782 1701
rect 1794 1698 1870 1701
rect 1906 1698 1998 1701
rect 2058 1698 2094 1701
rect 2122 1698 2134 1701
rect 2202 1698 2278 1701
rect 2282 1698 2350 1701
rect 2362 1698 2366 1701
rect 2386 1698 2486 1701
rect 2514 1698 2542 1701
rect 2554 1698 2574 1701
rect 2602 1698 2614 1701
rect 2746 1698 2782 1701
rect 2786 1698 2806 1701
rect 2810 1698 3025 1701
rect 3098 1698 3414 1701
rect 3474 1698 3486 1701
rect 798 1692 801 1698
rect 242 1688 278 1691
rect 322 1688 350 1691
rect 354 1688 598 1691
rect 602 1688 638 1691
rect 650 1688 782 1691
rect 818 1688 822 1691
rect 850 1688 902 1691
rect 926 1688 934 1691
rect 938 1688 966 1691
rect 982 1691 985 1698
rect 982 1688 1014 1691
rect 1042 1688 1294 1691
rect 1306 1688 1430 1691
rect 1526 1688 1598 1691
rect 1658 1688 1662 1691
rect 1682 1688 1702 1691
rect 1706 1688 1713 1691
rect 1722 1688 1798 1691
rect 1802 1688 1934 1691
rect 1954 1688 1974 1691
rect 1994 1688 2065 1691
rect 2090 1688 2126 1691
rect 2138 1688 2150 1691
rect 2158 1691 2161 1698
rect 2158 1688 2166 1691
rect 2230 1688 2238 1691
rect 2402 1688 2510 1691
rect 2546 1688 2550 1691
rect 2562 1688 2582 1691
rect 2594 1688 2625 1691
rect 114 1678 238 1681
rect 258 1678 270 1681
rect 330 1678 390 1681
rect 578 1678 630 1681
rect 662 1678 681 1681
rect 690 1678 694 1681
rect 714 1678 806 1681
rect 1058 1678 1062 1681
rect 1106 1678 1166 1681
rect 1202 1678 1326 1681
rect 1346 1678 1374 1681
rect 1526 1681 1529 1688
rect 2062 1682 2065 1688
rect 2230 1682 2233 1688
rect 2350 1682 2353 1688
rect 2622 1682 2625 1688
rect 2714 1688 2966 1691
rect 2978 1688 3006 1691
rect 3022 1691 3025 1698
rect 3526 1692 3529 1698
rect 3022 1688 3062 1691
rect 3162 1688 3166 1691
rect 3178 1688 3182 1691
rect 3210 1688 3214 1691
rect 3258 1688 3326 1691
rect 3330 1688 3358 1691
rect 3370 1688 3382 1691
rect 2686 1682 2689 1688
rect 1414 1678 1529 1681
rect 1554 1678 1638 1681
rect 1642 1678 1726 1681
rect 1746 1678 1822 1681
rect 1834 1678 1902 1681
rect 1906 1678 2006 1681
rect 2074 1678 2078 1681
rect 2106 1678 2214 1681
rect 2274 1678 2278 1681
rect 2322 1678 2334 1681
rect 2394 1678 2398 1681
rect 2410 1678 2414 1681
rect 2458 1678 2462 1681
rect 2546 1678 2590 1681
rect 2626 1678 2678 1681
rect 2714 1678 2718 1681
rect 2826 1678 2934 1681
rect 2978 1678 2982 1681
rect 3034 1678 3038 1681
rect 3166 1681 3169 1688
rect 3166 1678 3246 1681
rect 3266 1678 3310 1681
rect 3314 1678 3342 1681
rect 3354 1678 3358 1681
rect 3410 1678 3430 1681
rect 3454 1681 3457 1688
rect 3442 1678 3457 1681
rect 3502 1681 3505 1688
rect 3502 1678 3518 1681
rect 3522 1678 3526 1681
rect 3590 1681 3594 1682
rect 3562 1678 3594 1681
rect 42 1668 166 1671
rect 170 1668 182 1671
rect 226 1668 262 1671
rect 302 1671 305 1678
rect 298 1668 305 1671
rect 310 1672 313 1678
rect 662 1672 665 1678
rect 678 1672 681 1678
rect 1414 1672 1417 1678
rect 330 1668 358 1671
rect 426 1668 438 1671
rect 522 1668 529 1671
rect 538 1668 550 1671
rect 602 1668 638 1671
rect 806 1668 822 1671
rect 826 1668 846 1671
rect 850 1668 870 1671
rect 902 1668 926 1671
rect 970 1668 1030 1671
rect 1042 1668 1054 1671
rect 1090 1668 1150 1671
rect 1226 1668 1262 1671
rect 1266 1668 1318 1671
rect 1330 1668 1342 1671
rect 1358 1668 1366 1671
rect 1394 1668 1406 1671
rect 1450 1668 1462 1671
rect 1470 1668 1494 1671
rect 1522 1668 1702 1671
rect 1746 1668 1830 1671
rect 1850 1668 1854 1671
rect 1898 1668 1934 1671
rect 1946 1668 1966 1671
rect 1986 1668 2110 1671
rect 2158 1668 2182 1671
rect 2218 1668 2254 1671
rect 2274 1668 2470 1671
rect 2474 1668 2582 1671
rect 2586 1668 2614 1671
rect 2634 1668 2726 1671
rect 2730 1668 2782 1671
rect 2906 1668 2910 1671
rect 2938 1668 3254 1671
rect 3274 1668 3278 1671
rect 3298 1668 3374 1671
rect 3418 1668 3470 1671
rect 218 1658 222 1661
rect 258 1658 262 1661
rect 366 1661 369 1668
rect 526 1662 529 1668
rect 582 1662 585 1668
rect 806 1662 809 1668
rect 366 1658 414 1661
rect 418 1658 422 1661
rect 610 1658 614 1661
rect 626 1658 630 1661
rect 746 1658 750 1661
rect 770 1658 782 1661
rect 786 1658 798 1661
rect 834 1658 862 1661
rect 902 1661 905 1668
rect 1174 1662 1177 1668
rect 1214 1662 1217 1668
rect 1358 1662 1361 1668
rect 1430 1662 1433 1668
rect 1470 1662 1473 1668
rect 874 1658 905 1661
rect 914 1658 1094 1661
rect 1098 1658 1126 1661
rect 1186 1658 1198 1661
rect 1274 1658 1278 1661
rect 1338 1658 1342 1661
rect 1410 1658 1414 1661
rect 1438 1658 1454 1661
rect 1546 1658 1566 1661
rect 1602 1658 1606 1661
rect 1618 1658 1622 1661
rect 1674 1658 1678 1661
rect 1694 1658 1742 1661
rect 1754 1658 1766 1661
rect 1870 1661 1873 1668
rect 1850 1658 1873 1661
rect 1882 1658 1910 1661
rect 1930 1658 1934 1661
rect 1962 1658 1966 1661
rect 2158 1661 2161 1668
rect 1994 1658 2161 1661
rect 2170 1658 2174 1661
rect 2194 1658 2286 1661
rect 2290 1658 2465 1661
rect 2474 1658 2478 1661
rect 2498 1658 2518 1661
rect 2530 1658 2550 1661
rect 2578 1658 2582 1661
rect 2610 1658 2630 1661
rect 2662 1658 2750 1661
rect 2770 1658 2774 1661
rect 2802 1658 2814 1661
rect 2818 1658 2846 1661
rect 2882 1658 3030 1661
rect 3074 1658 3102 1661
rect 3106 1658 3142 1661
rect 3150 1658 3206 1661
rect 3378 1658 3398 1661
rect 3426 1658 3430 1661
rect 3434 1658 3454 1661
rect 158 1652 161 1658
rect 34 1648 110 1651
rect 186 1648 190 1651
rect 202 1648 222 1651
rect 338 1648 422 1651
rect 434 1648 446 1651
rect 454 1651 457 1658
rect 510 1652 513 1658
rect 1438 1652 1441 1658
rect 454 1648 486 1651
rect 514 1648 750 1651
rect 754 1648 774 1651
rect 834 1648 862 1651
rect 946 1648 1046 1651
rect 1258 1648 1278 1651
rect 1290 1648 1294 1651
rect 1318 1648 1326 1651
rect 1330 1648 1430 1651
rect 1538 1648 1558 1651
rect 1586 1648 1614 1651
rect 1638 1648 1646 1651
rect 1694 1651 1697 1658
rect 2182 1652 2185 1658
rect 2462 1652 2465 1658
rect 2654 1652 2657 1658
rect 2662 1652 2665 1658
rect 1650 1648 1697 1651
rect 1706 1648 1721 1651
rect 1730 1648 1822 1651
rect 1882 1648 1910 1651
rect 1946 1648 1958 1651
rect 1986 1648 1998 1651
rect 2050 1648 2078 1651
rect 2082 1648 2102 1651
rect 2122 1648 2126 1651
rect 2210 1648 2294 1651
rect 2306 1648 2398 1651
rect 2426 1648 2454 1651
rect 2466 1648 2641 1651
rect 2738 1648 2742 1651
rect 2894 1648 2926 1651
rect 2946 1648 2958 1651
rect 3058 1648 3086 1651
rect 3150 1651 3153 1658
rect 3138 1648 3153 1651
rect 3178 1648 3182 1651
rect 3194 1648 3310 1651
rect 3322 1648 3326 1651
rect 3366 1651 3369 1658
rect 3346 1648 3369 1651
rect 3394 1648 3398 1651
rect 3406 1648 3446 1651
rect 3474 1648 3494 1651
rect 182 1641 185 1648
rect 106 1638 185 1641
rect 206 1638 230 1641
rect 322 1638 342 1641
rect 538 1638 718 1641
rect 734 1638 846 1641
rect 890 1638 1134 1641
rect 1142 1638 1249 1641
rect 1258 1638 1710 1641
rect 1718 1641 1721 1648
rect 2110 1642 2113 1648
rect 2638 1642 2641 1648
rect 2894 1642 2897 1648
rect 3406 1642 3409 1648
rect 1718 1638 2054 1641
rect 2146 1638 2238 1641
rect 2274 1638 2326 1641
rect 2330 1638 2358 1641
rect 2362 1638 2574 1641
rect 2602 1638 2606 1641
rect 2682 1638 2830 1641
rect 2922 1638 3150 1641
rect 3182 1638 3198 1641
rect 3210 1638 3294 1641
rect 3362 1638 3382 1641
rect 206 1632 209 1638
rect 162 1628 166 1631
rect 726 1631 729 1638
rect 354 1628 729 1631
rect 734 1632 737 1638
rect 1142 1631 1145 1638
rect 786 1628 1145 1631
rect 1246 1631 1249 1638
rect 1246 1628 1350 1631
rect 1362 1628 1374 1631
rect 1386 1628 1390 1631
rect 1418 1628 1422 1631
rect 1442 1628 1454 1631
rect 1482 1628 1518 1631
rect 1522 1628 1534 1631
rect 1618 1628 1694 1631
rect 1710 1631 1713 1638
rect 1710 1628 2270 1631
rect 2282 1628 2302 1631
rect 2314 1628 2318 1631
rect 2338 1628 2342 1631
rect 2370 1628 2374 1631
rect 2426 1628 2438 1631
rect 2458 1628 2558 1631
rect 2570 1628 2774 1631
rect 2882 1628 2886 1631
rect 3182 1631 3185 1638
rect 2922 1628 3185 1631
rect 3490 1628 3518 1631
rect 170 1618 310 1621
rect 314 1618 398 1621
rect 758 1621 761 1628
rect 450 1618 609 1621
rect 758 1618 766 1621
rect 794 1618 1006 1621
rect 1026 1618 1126 1621
rect 154 1608 238 1611
rect 274 1608 278 1611
rect 394 1608 438 1611
rect 606 1611 609 1618
rect 1150 1612 1153 1628
rect 1178 1618 1254 1621
rect 1266 1618 1334 1621
rect 1362 1618 1374 1621
rect 1386 1618 1598 1621
rect 1610 1618 1718 1621
rect 1730 1618 1758 1621
rect 1818 1618 1870 1621
rect 1882 1618 1910 1621
rect 1922 1618 2142 1621
rect 2154 1618 2534 1621
rect 2642 1618 2718 1621
rect 2722 1618 3118 1621
rect 3190 1621 3193 1628
rect 3190 1618 3494 1621
rect 3134 1612 3137 1618
rect 606 1608 814 1611
rect 834 1608 846 1611
rect 850 1608 886 1611
rect 978 1608 1006 1611
rect 1010 1608 1046 1611
rect 1074 1608 1134 1611
rect 1242 1608 1254 1611
rect 1266 1608 1294 1611
rect 1402 1608 1502 1611
rect 1586 1608 1638 1611
rect 1682 1608 1702 1611
rect 1738 1608 1750 1611
rect 1770 1608 1774 1611
rect 1826 1608 1846 1611
rect 1850 1608 1894 1611
rect 1898 1608 2238 1611
rect 2242 1608 2422 1611
rect 2690 1608 2694 1611
rect 2730 1608 2750 1611
rect 2762 1608 3086 1611
rect 3194 1608 3198 1611
rect 3234 1608 3526 1611
rect 480 1603 482 1607
rect 486 1603 489 1607
rect 494 1603 496 1607
rect 542 1602 545 1608
rect 1512 1603 1514 1607
rect 1518 1603 1521 1607
rect 1526 1603 1528 1607
rect 2486 1602 2489 1608
rect 2536 1603 2538 1607
rect 2542 1603 2545 1607
rect 2550 1603 2552 1607
rect 194 1598 286 1601
rect 290 1598 294 1601
rect 314 1598 318 1601
rect 330 1598 334 1601
rect 386 1598 390 1601
rect 410 1598 470 1601
rect 562 1598 606 1601
rect 634 1598 638 1601
rect 682 1598 694 1601
rect 826 1598 1014 1601
rect 1018 1598 1110 1601
rect 1114 1598 1150 1601
rect 1154 1598 1174 1601
rect 1178 1598 1222 1601
rect 1250 1598 1350 1601
rect 1378 1598 1398 1601
rect 1434 1598 1494 1601
rect 1554 1598 1654 1601
rect 1674 1598 2326 1601
rect 2330 1598 2361 1601
rect 2650 1598 2694 1601
rect 2714 1598 2798 1601
rect 2826 1598 2990 1601
rect 3330 1598 3510 1601
rect 1366 1592 1369 1598
rect 2358 1592 2361 1598
rect 130 1588 534 1591
rect 538 1588 598 1591
rect 602 1588 854 1591
rect 858 1588 1038 1591
rect 1058 1588 1230 1591
rect 1234 1588 1262 1591
rect 1298 1588 1302 1591
rect 1322 1588 1334 1591
rect 1394 1588 1414 1591
rect 1434 1588 1470 1591
rect 1482 1588 2278 1591
rect 2302 1588 2310 1591
rect 2314 1588 2350 1591
rect 2370 1588 2422 1591
rect 2434 1588 2454 1591
rect 2466 1588 2494 1591
rect 2530 1588 2678 1591
rect 2802 1588 2857 1591
rect 2866 1588 2902 1591
rect 2978 1588 2998 1591
rect 3066 1588 3182 1591
rect 3186 1588 3350 1591
rect 3502 1588 3510 1591
rect 3514 1588 3558 1591
rect 2854 1582 2857 1588
rect 218 1578 662 1581
rect 674 1578 710 1581
rect 718 1578 726 1581
rect 730 1578 774 1581
rect 802 1578 918 1581
rect 930 1578 1078 1581
rect 1098 1578 1102 1581
rect 1122 1578 1278 1581
rect 1290 1578 1486 1581
rect 1506 1578 1566 1581
rect 1578 1578 1614 1581
rect 1626 1578 1630 1581
rect 1642 1578 1686 1581
rect 1714 1578 1726 1581
rect 1738 1578 1782 1581
rect 1802 1578 2134 1581
rect 2146 1578 2206 1581
rect 2226 1578 2254 1581
rect 2266 1578 2630 1581
rect 2978 1578 3337 1581
rect 3466 1578 3513 1581
rect 58 1568 150 1571
rect 194 1568 206 1571
rect 258 1568 286 1571
rect 290 1568 294 1571
rect 302 1568 310 1571
rect 314 1568 326 1571
rect 362 1568 374 1571
rect 418 1568 422 1571
rect 450 1568 462 1571
rect 474 1568 526 1571
rect 530 1568 534 1571
rect 570 1568 774 1571
rect 778 1568 838 1571
rect 866 1568 878 1571
rect 898 1568 910 1571
rect 926 1568 934 1571
rect 938 1568 982 1571
rect 1074 1568 1086 1571
rect 1138 1568 1142 1571
rect 1202 1568 1206 1571
rect 1226 1568 1230 1571
rect 1318 1568 1441 1571
rect 1450 1568 1478 1571
rect 1498 1568 1513 1571
rect 1522 1568 1590 1571
rect 1642 1568 1662 1571
rect 1706 1568 1886 1571
rect 1978 1568 2006 1571
rect 2014 1568 2022 1571
rect 2026 1568 2030 1571
rect 2058 1568 2142 1571
rect 2146 1568 2174 1571
rect 2186 1568 2214 1571
rect 2226 1568 2230 1571
rect 2242 1568 2382 1571
rect 2426 1568 2502 1571
rect 2514 1568 2542 1571
rect 2594 1568 2606 1571
rect 2738 1568 2742 1571
rect 2806 1571 2809 1578
rect 3334 1572 3337 1578
rect 3510 1572 3513 1578
rect 2806 1568 2838 1571
rect 2858 1568 2870 1571
rect 2946 1568 2990 1571
rect 3090 1568 3118 1571
rect 3154 1568 3158 1571
rect 3426 1568 3478 1571
rect 14 1561 17 1568
rect 398 1562 401 1568
rect 886 1562 889 1568
rect 14 1558 94 1561
rect 98 1558 102 1561
rect 138 1558 150 1561
rect 162 1558 198 1561
rect 266 1558 374 1561
rect 722 1558 726 1561
rect 802 1558 806 1561
rect 950 1558 1054 1561
rect 1318 1561 1321 1568
rect 1090 1558 1321 1561
rect 1338 1558 1342 1561
rect 1402 1558 1406 1561
rect 1426 1558 1430 1561
rect 1438 1561 1441 1568
rect 1438 1558 1462 1561
rect 1466 1558 1486 1561
rect 1490 1558 1502 1561
rect 1510 1561 1513 1568
rect 1894 1562 1897 1568
rect 1510 1558 1518 1561
rect 1522 1558 1534 1561
rect 1562 1558 1574 1561
rect 1594 1558 1606 1561
rect 1626 1558 1638 1561
rect 1650 1558 1702 1561
rect 1746 1558 1758 1561
rect 1802 1558 1830 1561
rect 1842 1558 1873 1561
rect 1882 1558 1886 1561
rect 1926 1558 2038 1561
rect 2066 1558 2097 1561
rect 2138 1558 2289 1561
rect 2298 1558 2302 1561
rect 2306 1558 2358 1561
rect 2418 1558 2422 1561
rect 2458 1558 2550 1561
rect 2562 1558 2582 1561
rect 2602 1558 2654 1561
rect 2666 1558 2734 1561
rect 2754 1558 2758 1561
rect 2878 1561 2881 1568
rect 2834 1558 2881 1561
rect 2894 1562 2897 1568
rect 2914 1558 2950 1561
rect 3074 1558 3078 1561
rect 3142 1561 3145 1568
rect 3142 1558 3166 1561
rect 3174 1561 3177 1568
rect 3174 1558 3278 1561
rect 3334 1561 3337 1568
rect 3334 1558 3366 1561
rect 3394 1558 3398 1561
rect 3402 1558 3478 1561
rect 118 1552 121 1558
rect 950 1552 953 1558
rect 1734 1552 1737 1558
rect 1766 1552 1769 1558
rect 42 1548 46 1551
rect 154 1548 214 1551
rect 226 1548 502 1551
rect 554 1548 574 1551
rect 586 1548 590 1551
rect 602 1548 630 1551
rect 658 1548 814 1551
rect 910 1548 918 1551
rect 922 1548 934 1551
rect 1034 1548 1046 1551
rect 1090 1548 1102 1551
rect 1210 1548 1217 1551
rect 1226 1548 1246 1551
rect 1266 1548 1318 1551
rect 1330 1548 1366 1551
rect 1450 1548 1470 1551
rect 1498 1548 1550 1551
rect 1578 1548 1582 1551
rect 1586 1548 1606 1551
rect 1610 1548 1686 1551
rect 1842 1548 1846 1551
rect 1870 1551 1873 1558
rect 1926 1551 1929 1558
rect 2054 1552 2057 1558
rect 2094 1552 2097 1558
rect 1870 1548 1929 1551
rect 1938 1548 1950 1551
rect 1970 1548 2022 1551
rect 2026 1548 2046 1551
rect 2126 1548 2134 1551
rect 2154 1548 2158 1551
rect 2194 1548 2262 1551
rect 2286 1551 2289 1558
rect 2286 1548 2366 1551
rect 2374 1551 2377 1558
rect 3550 1552 3553 1558
rect 2374 1548 2390 1551
rect 2450 1548 2454 1551
rect 2554 1548 2558 1551
rect 2570 1548 2574 1551
rect 2642 1548 2662 1551
rect 2714 1548 2846 1551
rect 2858 1548 2862 1551
rect 2874 1548 2878 1551
rect 2906 1548 3006 1551
rect 3066 1548 3070 1551
rect 3082 1548 3126 1551
rect 3130 1548 3230 1551
rect 3362 1548 3414 1551
rect 3418 1548 3534 1551
rect 3538 1548 3542 1551
rect 3590 1551 3594 1552
rect 3562 1548 3594 1551
rect 870 1542 873 1548
rect 26 1538 30 1541
rect 58 1538 198 1541
rect 322 1538 374 1541
rect 418 1538 446 1541
rect 490 1538 502 1541
rect 530 1538 534 1541
rect 538 1538 622 1541
rect 626 1538 654 1541
rect 698 1538 710 1541
rect 722 1538 742 1541
rect 754 1538 822 1541
rect 890 1538 942 1541
rect 986 1538 1022 1541
rect 1050 1538 1054 1541
rect 1066 1538 1094 1541
rect 1214 1541 1217 1548
rect 1694 1542 1697 1548
rect 1214 1538 1230 1541
rect 1306 1538 1334 1541
rect 1354 1538 1382 1541
rect 1410 1538 1414 1541
rect 1426 1538 1478 1541
rect 1490 1538 1502 1541
rect 1530 1538 1601 1541
rect 1610 1538 1614 1541
rect 1718 1541 1721 1548
rect 1718 1538 2094 1541
rect 2110 1541 2113 1548
rect 2106 1538 2113 1541
rect 2126 1542 2129 1548
rect 2598 1542 2601 1548
rect 2154 1538 2190 1541
rect 2266 1538 2310 1541
rect 2362 1538 2382 1541
rect 2402 1538 2414 1541
rect 2450 1538 2574 1541
rect 2602 1538 2686 1541
rect 2734 1538 2934 1541
rect 2946 1538 2990 1541
rect 3138 1538 3222 1541
rect 3226 1538 3233 1541
rect 3346 1538 3438 1541
rect 3466 1538 3470 1541
rect 286 1532 289 1538
rect 154 1528 158 1531
rect 178 1528 190 1531
rect 298 1528 358 1531
rect 370 1528 377 1531
rect 486 1531 489 1538
rect 426 1528 489 1531
rect 578 1528 582 1531
rect 610 1528 614 1531
rect 822 1531 825 1538
rect 626 1528 769 1531
rect 822 1528 870 1531
rect 874 1528 910 1531
rect 930 1528 934 1531
rect 962 1528 1142 1531
rect 1154 1528 1158 1531
rect 1178 1528 1182 1531
rect 1250 1528 1254 1531
rect 1298 1528 1310 1531
rect 1346 1528 1350 1531
rect 1402 1528 1422 1531
rect 1426 1528 1454 1531
rect 1482 1528 1526 1531
rect 1546 1528 1550 1531
rect 1598 1531 1601 1538
rect 1630 1532 1633 1538
rect 1678 1532 1681 1538
rect 1598 1528 1625 1531
rect 1690 1528 1769 1531
rect 1778 1528 1806 1531
rect 1810 1528 1862 1531
rect 1898 1528 1918 1531
rect 1938 1528 1942 1531
rect 1986 1528 1990 1531
rect 2026 1528 2038 1531
rect 2090 1528 2110 1531
rect 2218 1528 2222 1531
rect 2242 1528 2246 1531
rect 2266 1528 2278 1531
rect 2290 1528 2294 1531
rect 2346 1528 2406 1531
rect 2410 1528 2526 1531
rect 2582 1531 2585 1538
rect 2734 1532 2737 1538
rect 2546 1528 2585 1531
rect 2602 1528 2622 1531
rect 2642 1528 2646 1531
rect 2762 1528 2790 1531
rect 2818 1528 2822 1531
rect 2866 1528 2894 1531
rect 2898 1528 2910 1531
rect 3070 1531 3073 1538
rect 2938 1528 3073 1531
rect 3146 1528 3150 1531
rect 3178 1528 3214 1531
rect 3346 1528 3478 1531
rect 3498 1528 3502 1531
rect 374 1522 377 1528
rect 170 1518 174 1521
rect 250 1518 342 1521
rect 402 1518 446 1521
rect 506 1518 686 1521
rect 702 1518 710 1521
rect 714 1518 750 1521
rect 766 1521 769 1528
rect 1262 1522 1265 1528
rect 1286 1522 1289 1528
rect 766 1518 958 1521
rect 1090 1518 1126 1521
rect 1138 1518 1150 1521
rect 1178 1518 1206 1521
rect 1306 1518 1382 1521
rect 1402 1518 1430 1521
rect 1482 1518 1542 1521
rect 1554 1518 1558 1521
rect 1586 1518 1614 1521
rect 1622 1521 1625 1528
rect 1766 1522 1769 1528
rect 2454 1522 2457 1528
rect 1622 1518 1638 1521
rect 1642 1518 1654 1521
rect 1690 1518 1758 1521
rect 1778 1518 1790 1521
rect 1826 1518 1862 1521
rect 1890 1518 1910 1521
rect 1946 1518 1990 1521
rect 2010 1518 2105 1521
rect 2114 1518 2446 1521
rect 2514 1518 2518 1521
rect 2578 1518 2662 1521
rect 2670 1521 2673 1528
rect 2734 1522 2737 1528
rect 2806 1522 2809 1528
rect 2926 1522 2929 1528
rect 2670 1518 2726 1521
rect 2946 1518 2974 1521
rect 2978 1518 2998 1521
rect 3002 1518 3030 1521
rect 3102 1521 3105 1528
rect 3034 1518 3105 1521
rect 3186 1518 3230 1521
rect 3338 1518 3350 1521
rect 3426 1518 3430 1521
rect 1022 1512 1025 1518
rect 114 1508 310 1511
rect 330 1508 334 1511
rect 354 1508 630 1511
rect 642 1508 694 1511
rect 746 1508 758 1511
rect 858 1508 862 1511
rect 882 1508 918 1511
rect 930 1508 982 1511
rect 1034 1508 1166 1511
rect 1462 1511 1465 1518
rect 1202 1508 1465 1511
rect 1482 1508 1494 1511
rect 1498 1508 1566 1511
rect 1578 1508 1646 1511
rect 1674 1508 1686 1511
rect 1698 1508 1758 1511
rect 1770 1508 1790 1511
rect 1798 1508 1830 1511
rect 1842 1508 1846 1511
rect 1858 1508 1870 1511
rect 1882 1508 1950 1511
rect 1954 1508 1974 1511
rect 1994 1508 2014 1511
rect 2082 1508 2086 1511
rect 2102 1511 2105 1518
rect 3382 1512 3385 1518
rect 2102 1508 2134 1511
rect 2138 1508 2150 1511
rect 2162 1508 2486 1511
rect 2490 1508 2718 1511
rect 2762 1508 2854 1511
rect 2922 1508 2926 1511
rect 2938 1508 2950 1511
rect 3130 1508 3206 1511
rect 3274 1508 3302 1511
rect 3466 1508 3470 1511
rect 992 1503 994 1507
rect 998 1503 1001 1507
rect 1006 1503 1008 1507
rect 1662 1502 1665 1508
rect 258 1498 350 1501
rect 362 1498 582 1501
rect 642 1498 646 1501
rect 770 1498 822 1501
rect 842 1498 982 1501
rect 1106 1498 1118 1501
rect 1138 1498 1246 1501
rect 1258 1498 1270 1501
rect 1298 1498 1342 1501
rect 1354 1498 1446 1501
rect 1454 1498 1614 1501
rect 1626 1498 1646 1501
rect 1798 1501 1801 1508
rect 2024 1503 2026 1507
rect 2030 1503 2033 1507
rect 2038 1503 2040 1507
rect 3040 1503 3042 1507
rect 3046 1503 3049 1507
rect 3054 1503 3056 1507
rect 3446 1502 3449 1508
rect 1730 1498 1801 1501
rect 1826 1498 1886 1501
rect 1914 1498 2014 1501
rect 2098 1498 2102 1501
rect 2122 1498 2166 1501
rect 2170 1498 2230 1501
rect 2234 1498 2310 1501
rect 2354 1498 2366 1501
rect 2482 1498 2534 1501
rect 2562 1498 2582 1501
rect 2594 1498 2638 1501
rect 2642 1498 2678 1501
rect 2730 1498 2734 1501
rect 2794 1498 2950 1501
rect 3002 1498 3022 1501
rect 3234 1498 3398 1501
rect 82 1488 390 1491
rect 394 1488 438 1491
rect 446 1488 454 1491
rect 702 1488 822 1491
rect 1034 1488 1134 1491
rect 1194 1488 1198 1491
rect 1214 1488 1222 1491
rect 1226 1488 1302 1491
rect 1322 1488 1385 1491
rect 1394 1488 1414 1491
rect 1454 1491 1457 1498
rect 1426 1488 1457 1491
rect 1466 1488 1625 1491
rect 1630 1488 1638 1491
rect 1650 1488 1694 1491
rect 1714 1488 1734 1491
rect 1762 1488 1774 1491
rect 1786 1488 1798 1491
rect 1810 1488 1822 1491
rect 2118 1491 2121 1498
rect 1842 1488 2121 1491
rect 2194 1488 2198 1491
rect 2210 1488 2286 1491
rect 2314 1488 2334 1491
rect 2362 1488 2630 1491
rect 2666 1488 2686 1491
rect 2890 1488 2902 1491
rect 2906 1488 2942 1491
rect 2994 1488 3142 1491
rect 3170 1488 3486 1491
rect 702 1482 705 1488
rect 178 1478 206 1481
rect 210 1478 214 1481
rect 346 1478 374 1481
rect 418 1478 422 1481
rect 602 1478 654 1481
rect 754 1478 838 1481
rect 886 1481 889 1488
rect 886 1478 894 1481
rect 922 1478 942 1481
rect 954 1478 974 1481
rect 986 1478 1030 1481
rect 1066 1478 1070 1481
rect 1074 1478 1166 1481
rect 1242 1478 1262 1481
rect 1270 1478 1278 1481
rect 1282 1478 1302 1481
rect 1306 1478 1334 1481
rect 1346 1478 1358 1481
rect 1382 1481 1385 1488
rect 1382 1478 1398 1481
rect 1418 1478 1446 1481
rect 1458 1478 1574 1481
rect 1622 1481 1625 1488
rect 2358 1482 2361 1488
rect 1622 1478 1678 1481
rect 1706 1478 1726 1481
rect 1730 1478 1742 1481
rect 1786 1478 1790 1481
rect 1818 1478 1902 1481
rect 1930 1478 1966 1481
rect 1994 1478 1998 1481
rect 2010 1478 2134 1481
rect 2218 1478 2230 1481
rect 2274 1478 2278 1481
rect 2286 1478 2334 1481
rect 2370 1478 2406 1481
rect 2410 1478 2462 1481
rect 2482 1478 2494 1481
rect 2498 1478 2582 1481
rect 2606 1478 2670 1481
rect 2726 1481 2729 1488
rect 2822 1481 2825 1488
rect 2726 1478 2825 1481
rect 2850 1478 2862 1481
rect 2882 1478 2886 1481
rect 2906 1478 2966 1481
rect 2978 1478 3006 1481
rect 3010 1478 3017 1481
rect 3026 1478 3166 1481
rect 3270 1478 3278 1481
rect 3282 1478 3286 1481
rect 3298 1478 3366 1481
rect 3370 1478 3374 1481
rect 3402 1478 3422 1481
rect 3442 1478 3454 1481
rect 3458 1478 3502 1481
rect 3514 1478 3542 1481
rect 58 1468 94 1471
rect 202 1468 302 1471
rect 306 1468 414 1471
rect 426 1468 462 1471
rect 498 1468 558 1471
rect 562 1468 598 1471
rect 618 1468 646 1471
rect 714 1468 734 1471
rect 770 1468 814 1471
rect 910 1471 913 1478
rect 2286 1472 2289 1478
rect 2606 1472 2609 1478
rect 874 1468 913 1471
rect 958 1468 1022 1471
rect 1058 1468 1174 1471
rect 1178 1468 1214 1471
rect 1242 1468 1286 1471
rect 1294 1468 1454 1471
rect 1458 1468 1486 1471
rect 1506 1468 1510 1471
rect 1546 1468 1582 1471
rect 1610 1468 1614 1471
rect 1634 1468 1710 1471
rect 1730 1468 1758 1471
rect 1770 1468 1854 1471
rect 1866 1468 1870 1471
rect 1874 1468 2046 1471
rect 2054 1468 2097 1471
rect 2106 1468 2118 1471
rect 2178 1468 2182 1471
rect 2258 1468 2286 1471
rect 2362 1468 2425 1471
rect 2434 1468 2558 1471
rect 2586 1468 2606 1471
rect 2666 1468 2678 1471
rect 2738 1468 2742 1471
rect 2762 1468 2798 1471
rect 2822 1468 2865 1471
rect 2874 1468 2894 1471
rect 2954 1468 2982 1471
rect 2986 1468 3030 1471
rect 3058 1468 3070 1471
rect 3234 1468 3334 1471
rect 3338 1468 3374 1471
rect 3402 1468 3406 1471
rect 3510 1471 3513 1478
rect 3418 1468 3513 1471
rect 3522 1468 3526 1471
rect 926 1462 929 1468
rect 82 1458 94 1461
rect 138 1458 190 1461
rect 266 1458 286 1461
rect 298 1458 326 1461
rect 362 1458 414 1461
rect 418 1458 446 1461
rect 522 1458 534 1461
rect 538 1458 558 1461
rect 602 1458 662 1461
rect 698 1458 830 1461
rect 834 1458 902 1461
rect 906 1458 926 1461
rect 958 1461 961 1468
rect 930 1458 961 1461
rect 970 1458 998 1461
rect 1010 1458 1022 1461
rect 1058 1458 1126 1461
rect 1138 1458 1158 1461
rect 1162 1458 1166 1461
rect 1186 1458 1222 1461
rect 1294 1461 1297 1468
rect 1282 1458 1297 1461
rect 1306 1458 1310 1461
rect 1370 1458 1382 1461
rect 1406 1458 1433 1461
rect 1450 1458 1462 1461
rect 1474 1458 1534 1461
rect 1570 1458 1582 1461
rect 1594 1458 1622 1461
rect 1642 1458 1726 1461
rect 1746 1458 1758 1461
rect 1770 1458 1822 1461
rect 1834 1458 1902 1461
rect 1910 1458 1918 1461
rect 1922 1458 1998 1461
rect 2054 1461 2057 1468
rect 2002 1458 2057 1461
rect 2074 1458 2078 1461
rect 2094 1461 2097 1468
rect 2094 1458 2110 1461
rect 2114 1458 2126 1461
rect 2150 1461 2153 1468
rect 2422 1462 2425 1468
rect 2150 1458 2190 1461
rect 2202 1458 2206 1461
rect 2210 1458 2214 1461
rect 2250 1458 2270 1461
rect 2282 1458 2318 1461
rect 2338 1458 2406 1461
rect 2454 1458 2510 1461
rect 2514 1458 2550 1461
rect 2562 1458 2598 1461
rect 2682 1458 2686 1461
rect 2710 1461 2713 1468
rect 2690 1458 2713 1461
rect 2762 1458 2774 1461
rect 2822 1461 2825 1468
rect 2778 1458 2825 1461
rect 2834 1458 2846 1461
rect 2862 1461 2865 1468
rect 2862 1458 2886 1461
rect 2910 1461 2913 1468
rect 2898 1458 2913 1461
rect 2926 1462 2929 1468
rect 2966 1458 2974 1461
rect 2978 1459 3110 1461
rect 2978 1458 3113 1459
rect 3186 1458 3206 1461
rect 3226 1458 3238 1461
rect 3250 1458 3254 1461
rect 3266 1458 3294 1461
rect 3322 1458 3494 1461
rect 254 1452 257 1458
rect 1198 1452 1201 1458
rect 106 1448 110 1451
rect 146 1448 150 1451
rect 162 1448 166 1451
rect 258 1448 318 1451
rect 330 1448 390 1451
rect 402 1448 430 1451
rect 434 1448 550 1451
rect 554 1448 598 1451
rect 610 1448 638 1451
rect 762 1448 766 1451
rect 802 1448 830 1451
rect 834 1448 926 1451
rect 994 1448 1030 1451
rect 1074 1448 1086 1451
rect 1098 1448 1126 1451
rect 1246 1451 1249 1458
rect 1262 1451 1265 1458
rect 1246 1448 1265 1451
rect 1406 1451 1409 1458
rect 1430 1452 1433 1458
rect 2142 1452 2145 1458
rect 2454 1452 2457 1458
rect 1274 1448 1409 1451
rect 1418 1448 1425 1451
rect 1458 1448 1462 1451
rect 1482 1448 1542 1451
rect 1554 1448 1590 1451
rect 1594 1448 1606 1451
rect 1634 1448 1646 1451
rect 1674 1448 1702 1451
rect 1714 1448 1718 1451
rect 1738 1448 1750 1451
rect 1770 1448 2006 1451
rect 2034 1448 2094 1451
rect 2122 1448 2126 1451
rect 2178 1448 2198 1451
rect 2202 1448 2206 1451
rect 2386 1448 2414 1451
rect 2426 1448 2430 1451
rect 2470 1448 2542 1451
rect 2570 1448 2670 1451
rect 2690 1448 2718 1451
rect 2770 1448 2774 1451
rect 2890 1448 2958 1451
rect 2970 1448 3030 1451
rect 3066 1448 3166 1451
rect 3218 1448 3230 1451
rect 3234 1448 3414 1451
rect 3418 1448 3422 1451
rect 3474 1448 3558 1451
rect 3590 1451 3594 1452
rect 3562 1448 3594 1451
rect 98 1438 126 1441
rect 170 1438 222 1441
rect 234 1438 390 1441
rect 418 1438 478 1441
rect 538 1438 590 1441
rect 594 1438 622 1441
rect 650 1438 718 1441
rect 746 1438 774 1441
rect 826 1438 878 1441
rect 930 1438 1006 1441
rect 1066 1438 1158 1441
rect 1234 1438 1278 1441
rect 1290 1438 1342 1441
rect 1386 1438 1414 1441
rect 1422 1441 1425 1448
rect 1422 1438 1486 1441
rect 1498 1438 1502 1441
rect 1562 1438 1614 1441
rect 1670 1441 1673 1448
rect 1726 1442 1729 1448
rect 1618 1438 1673 1441
rect 1682 1438 1694 1441
rect 1754 1438 1918 1441
rect 1930 1438 1934 1441
rect 1962 1438 1990 1441
rect 1994 1438 2086 1441
rect 2254 1441 2257 1448
rect 2470 1442 2473 1448
rect 2090 1438 2294 1441
rect 2306 1438 2366 1441
rect 2482 1438 2558 1441
rect 2794 1438 3062 1441
rect 3154 1438 3190 1441
rect 3274 1438 3318 1441
rect 3354 1438 3358 1441
rect 3434 1438 3550 1441
rect 62 1431 65 1438
rect 62 1428 326 1431
rect 354 1428 398 1431
rect 450 1428 454 1431
rect 478 1428 726 1431
rect 782 1431 785 1438
rect 1022 1432 1025 1438
rect 782 1428 838 1431
rect 978 1428 1006 1431
rect 1082 1428 1110 1431
rect 1174 1431 1177 1438
rect 1174 1428 1542 1431
rect 1546 1428 1774 1431
rect 1786 1428 1798 1431
rect 1802 1428 1854 1431
rect 1858 1428 1878 1431
rect 1882 1428 1958 1431
rect 2002 1428 2030 1431
rect 2074 1428 2078 1431
rect 2098 1428 2238 1431
rect 2250 1428 2934 1431
rect 3190 1431 3193 1438
rect 3190 1428 3246 1431
rect 3250 1428 3366 1431
rect 478 1421 481 1428
rect 1118 1422 1121 1428
rect 2990 1422 2993 1428
rect 314 1418 481 1421
rect 514 1418 942 1421
rect 1034 1418 1086 1421
rect 1154 1418 1190 1421
rect 1210 1418 1254 1421
rect 1274 1418 1294 1421
rect 1330 1418 1350 1421
rect 1362 1418 1406 1421
rect 1418 1418 1422 1421
rect 1502 1418 1590 1421
rect 1602 1418 1694 1421
rect 1714 1418 1734 1421
rect 1746 1418 1774 1421
rect 1810 1418 1838 1421
rect 1850 1418 1966 1421
rect 1970 1418 2814 1421
rect 2866 1418 2910 1421
rect 3054 1421 3057 1428
rect 3054 1418 3286 1421
rect 3290 1418 3342 1421
rect 3346 1418 3358 1421
rect 3366 1421 3369 1428
rect 3366 1418 3382 1421
rect 3458 1418 3542 1421
rect 266 1408 318 1411
rect 1502 1411 1505 1418
rect 586 1408 1505 1411
rect 1538 1408 1849 1411
rect 480 1403 482 1407
rect 486 1403 489 1407
rect 494 1403 496 1407
rect 1512 1403 1514 1407
rect 1518 1403 1521 1407
rect 1526 1403 1528 1407
rect 1846 1402 1849 1408
rect 1922 1408 1934 1411
rect 1946 1408 1950 1411
rect 1954 1408 1998 1411
rect 2010 1408 2102 1411
rect 2114 1408 2246 1411
rect 2258 1408 2406 1411
rect 2418 1408 2470 1411
rect 2474 1408 2510 1411
rect 2562 1408 2590 1411
rect 2634 1408 2910 1411
rect 3434 1408 3454 1411
rect 3466 1408 3542 1411
rect 1870 1402 1873 1408
rect 2536 1403 2538 1407
rect 2542 1403 2545 1407
rect 2550 1403 2552 1407
rect 282 1398 398 1401
rect 562 1398 750 1401
rect 794 1398 958 1401
rect 1002 1398 1014 1401
rect 1026 1398 1270 1401
rect 1282 1398 1302 1401
rect 1314 1398 1502 1401
rect 1586 1398 1646 1401
rect 1650 1398 1694 1401
rect 1714 1398 1718 1401
rect 1746 1398 1750 1401
rect 1786 1398 1806 1401
rect 1922 1398 1966 1401
rect 2058 1398 2086 1401
rect 2142 1398 2166 1401
rect 2178 1398 2238 1401
rect 2282 1398 2310 1401
rect 2370 1398 2382 1401
rect 2450 1398 2510 1401
rect 2642 1398 2694 1401
rect 2698 1398 2862 1401
rect 3106 1398 3342 1401
rect 3346 1398 3390 1401
rect 234 1388 246 1391
rect 314 1388 494 1391
rect 642 1388 782 1391
rect 810 1388 870 1391
rect 894 1388 969 1391
rect 978 1388 1078 1391
rect 1130 1388 1158 1391
rect 1170 1388 1174 1391
rect 1250 1388 1681 1391
rect 1690 1388 1798 1391
rect 1818 1388 2070 1391
rect 2142 1391 2145 1398
rect 2082 1388 2145 1391
rect 2154 1388 2158 1391
rect 2170 1388 2174 1391
rect 2178 1388 2182 1391
rect 2194 1388 2222 1391
rect 2278 1391 2281 1398
rect 2234 1388 2281 1391
rect 2298 1388 2350 1391
rect 2410 1388 2502 1391
rect 2578 1388 2614 1391
rect 2674 1388 2702 1391
rect 2730 1388 2838 1391
rect 2866 1388 3206 1391
rect 3210 1388 3278 1391
rect 3338 1388 3406 1391
rect 894 1382 897 1388
rect 242 1378 342 1381
rect 346 1378 358 1381
rect 378 1378 486 1381
rect 658 1378 798 1381
rect 802 1378 870 1381
rect 914 1378 958 1381
rect 966 1381 969 1388
rect 966 1378 1022 1381
rect 1042 1378 1062 1381
rect 1090 1378 1230 1381
rect 1242 1378 1262 1381
rect 1266 1378 1430 1381
rect 1434 1378 1558 1381
rect 1578 1378 1638 1381
rect 1650 1378 1654 1381
rect 1678 1381 1681 1388
rect 1678 1378 1822 1381
rect 1850 1378 1902 1381
rect 1914 1378 2014 1381
rect 2018 1378 2102 1381
rect 2210 1378 2342 1381
rect 2354 1378 2825 1381
rect 2834 1378 2886 1381
rect 2890 1378 2897 1381
rect 2906 1378 2998 1381
rect 3234 1378 3470 1381
rect 3486 1378 3534 1381
rect 238 1372 241 1378
rect 58 1368 70 1371
rect 106 1368 142 1371
rect 170 1368 182 1371
rect 306 1368 318 1371
rect 450 1368 526 1371
rect 606 1371 609 1378
rect 606 1368 782 1371
rect 786 1368 798 1371
rect 802 1368 838 1371
rect 858 1368 878 1371
rect 898 1368 942 1371
rect 970 1368 1190 1371
rect 1226 1368 1662 1371
rect 1674 1368 1766 1371
rect 1834 1368 1886 1371
rect 1914 1368 1942 1371
rect 1954 1368 1974 1371
rect 2034 1368 2046 1371
rect 2090 1368 2102 1371
rect 2146 1368 2198 1371
rect 2258 1368 2374 1371
rect 2394 1368 2518 1371
rect 2530 1368 2625 1371
rect 42 1358 110 1361
rect 114 1358 310 1361
rect 362 1358 366 1361
rect 422 1361 425 1368
rect 566 1362 569 1368
rect 394 1358 425 1361
rect 442 1358 462 1361
rect 538 1358 558 1361
rect 570 1358 606 1361
rect 698 1358 926 1361
rect 970 1358 990 1361
rect 1002 1358 1062 1361
rect 1066 1358 1134 1361
rect 1162 1358 1262 1361
rect 1274 1358 1286 1361
rect 1306 1358 1342 1361
rect 1370 1358 1454 1361
rect 1498 1358 1505 1361
rect 1522 1358 1574 1361
rect 1610 1358 1705 1361
rect 1714 1358 1726 1361
rect 1822 1361 1825 1368
rect 1894 1362 1897 1368
rect 2622 1362 2625 1368
rect 2742 1368 2782 1371
rect 2822 1371 2825 1378
rect 2822 1368 3030 1371
rect 3034 1368 3134 1371
rect 3486 1371 3489 1378
rect 3274 1368 3489 1371
rect 3494 1368 3502 1371
rect 3506 1368 3526 1371
rect 1818 1358 1825 1361
rect 1874 1358 1878 1361
rect 1902 1358 1910 1361
rect 1974 1358 2014 1361
rect 2050 1358 2110 1361
rect 2186 1358 2190 1361
rect 2202 1358 2230 1361
rect 2362 1358 2366 1361
rect 2370 1358 2478 1361
rect 2498 1358 2502 1361
rect 2530 1358 2542 1361
rect 2594 1358 2598 1361
rect 2726 1361 2729 1368
rect 2706 1358 2729 1361
rect 2742 1362 2745 1368
rect 2762 1358 2766 1361
rect 2794 1358 2838 1361
rect 2930 1358 2942 1361
rect 2986 1358 3086 1361
rect 3094 1358 3190 1361
rect 3194 1358 3286 1361
rect 3338 1358 3478 1361
rect 3482 1358 3510 1361
rect 686 1352 689 1358
rect 50 1348 70 1351
rect 74 1348 142 1351
rect 146 1348 166 1351
rect 170 1348 190 1351
rect 258 1348 318 1351
rect 370 1348 446 1351
rect 458 1348 462 1351
rect 506 1348 537 1351
rect 706 1348 726 1351
rect 730 1348 737 1351
rect 762 1348 846 1351
rect 850 1348 902 1351
rect 978 1348 1006 1351
rect 1018 1348 1073 1351
rect 1098 1348 1118 1351
rect 1186 1348 1206 1351
rect 1218 1348 1238 1351
rect 1242 1348 1326 1351
rect 1358 1351 1361 1358
rect 1502 1352 1505 1358
rect 1598 1352 1601 1358
rect 1346 1348 1374 1351
rect 1386 1348 1390 1351
rect 1402 1348 1438 1351
rect 1530 1348 1534 1351
rect 1578 1348 1582 1351
rect 1634 1348 1646 1351
rect 1690 1348 1694 1351
rect 1702 1351 1705 1358
rect 1902 1352 1905 1358
rect 1918 1352 1921 1358
rect 1942 1352 1945 1358
rect 1974 1352 1977 1358
rect 2614 1352 2617 1358
rect 2686 1352 2689 1358
rect 1702 1348 1734 1351
rect 1762 1348 1766 1351
rect 1778 1348 1782 1351
rect 1786 1348 1886 1351
rect 2058 1348 2062 1351
rect 2098 1348 2102 1351
rect 2218 1348 2254 1351
rect 2266 1348 2270 1351
rect 2330 1348 2342 1351
rect 2394 1348 2398 1351
rect 2402 1348 2406 1351
rect 2426 1348 2430 1351
rect 2506 1348 2510 1351
rect 2578 1348 2582 1351
rect 2762 1348 2814 1351
rect 2826 1348 2830 1351
rect 2858 1348 2862 1351
rect 2954 1348 2958 1351
rect 2962 1348 2982 1351
rect 3002 1348 3006 1351
rect 3094 1351 3097 1358
rect 3078 1348 3097 1351
rect 3138 1348 3166 1351
rect 3170 1348 3230 1351
rect 3234 1348 3454 1351
rect 3590 1351 3594 1352
rect 3458 1348 3594 1351
rect 534 1342 537 1348
rect 910 1342 913 1348
rect 34 1338 94 1341
rect 98 1338 126 1341
rect 238 1338 254 1341
rect 330 1338 342 1341
rect 442 1338 454 1341
rect 562 1338 582 1341
rect 586 1338 622 1341
rect 626 1338 718 1341
rect 826 1338 862 1341
rect 946 1338 950 1341
rect 986 1338 1006 1341
rect 1026 1338 1038 1341
rect 1070 1341 1073 1348
rect 1982 1342 1985 1348
rect 1070 1338 1086 1341
rect 1146 1338 1150 1341
rect 1154 1338 1310 1341
rect 1330 1338 1342 1341
rect 1354 1338 1718 1341
rect 1762 1338 1766 1341
rect 1834 1338 1966 1341
rect 2042 1338 2113 1341
rect 2122 1338 2270 1341
rect 2314 1338 2510 1341
rect 2530 1338 2577 1341
rect 238 1331 241 1338
rect 114 1328 241 1331
rect 250 1328 262 1331
rect 310 1331 313 1338
rect 1990 1332 1993 1338
rect 2110 1332 2113 1338
rect 2574 1332 2577 1338
rect 2602 1338 2638 1341
rect 2658 1338 2678 1341
rect 2726 1341 2729 1348
rect 3078 1342 3081 1348
rect 3454 1342 3457 1348
rect 2706 1338 2729 1341
rect 2738 1338 2742 1341
rect 2754 1338 2758 1341
rect 2802 1338 2806 1341
rect 2818 1338 2926 1341
rect 2930 1338 2966 1341
rect 2970 1338 3006 1341
rect 3114 1338 3230 1341
rect 3234 1338 3238 1341
rect 3274 1338 3278 1341
rect 3338 1338 3350 1341
rect 3362 1338 3377 1341
rect 2582 1332 2585 1338
rect 3086 1332 3089 1338
rect 3374 1332 3377 1338
rect 3434 1338 3438 1341
rect 3474 1338 3494 1341
rect 3538 1338 3542 1341
rect 3406 1332 3409 1338
rect 310 1328 358 1331
rect 378 1328 438 1331
rect 602 1328 742 1331
rect 834 1328 838 1331
rect 842 1328 878 1331
rect 954 1328 1030 1331
rect 1050 1328 1054 1331
rect 1106 1328 1150 1331
rect 1162 1328 1182 1331
rect 1210 1328 1214 1331
rect 1226 1328 1334 1331
rect 1362 1328 1366 1331
rect 1386 1328 1398 1331
rect 1442 1328 1470 1331
rect 1570 1328 1574 1331
rect 1634 1328 1678 1331
rect 1690 1328 1694 1331
rect 1730 1328 1734 1331
rect 1762 1328 1830 1331
rect 1838 1328 1846 1331
rect 1878 1328 1886 1331
rect 1890 1328 1918 1331
rect 1938 1328 1950 1331
rect 2066 1328 2078 1331
rect 2098 1328 2102 1331
rect 2190 1328 2198 1331
rect 2202 1328 2214 1331
rect 2226 1328 2294 1331
rect 2306 1328 2358 1331
rect 2370 1328 2382 1331
rect 2386 1328 2470 1331
rect 2506 1328 2566 1331
rect 2602 1328 2622 1331
rect 2678 1328 2686 1331
rect 2690 1328 2694 1331
rect 2714 1328 2766 1331
rect 2802 1328 2822 1331
rect 2842 1328 2918 1331
rect 2926 1328 2958 1331
rect 3002 1328 3070 1331
rect 3178 1328 3246 1331
rect 3306 1328 3310 1331
rect 3354 1328 3358 1331
rect 3426 1328 3470 1331
rect 3482 1328 3486 1331
rect 3490 1328 3502 1331
rect 258 1318 350 1321
rect 450 1318 646 1321
rect 666 1318 742 1321
rect 866 1318 1049 1321
rect 1198 1321 1201 1328
rect 1406 1322 1409 1328
rect 1082 1318 1193 1321
rect 1198 1318 1270 1321
rect 1282 1318 1342 1321
rect 1354 1318 1390 1321
rect 1418 1318 1518 1321
rect 1562 1318 1606 1321
rect 1646 1318 1654 1321
rect 1658 1318 1694 1321
rect 1706 1318 1806 1321
rect 1826 1318 1926 1321
rect 1938 1318 1942 1321
rect 1994 1318 2030 1321
rect 2038 1321 2041 1328
rect 2126 1322 2129 1328
rect 2166 1322 2169 1328
rect 2654 1322 2657 1328
rect 2926 1322 2929 1328
rect 2038 1318 2046 1321
rect 2074 1318 2078 1321
rect 2082 1318 2118 1321
rect 2226 1318 2230 1321
rect 2242 1318 2246 1321
rect 2490 1318 2494 1321
rect 2514 1318 2646 1321
rect 2706 1318 2718 1321
rect 2850 1318 2854 1321
rect 2974 1321 2977 1328
rect 2946 1318 2977 1321
rect 2994 1318 3198 1321
rect 3202 1318 3206 1321
rect 3218 1318 3310 1321
rect 3354 1318 3462 1321
rect 66 1308 526 1311
rect 554 1308 662 1311
rect 706 1308 846 1311
rect 882 1308 982 1311
rect 1046 1311 1049 1318
rect 1046 1308 1102 1311
rect 1138 1308 1174 1311
rect 1190 1311 1193 1318
rect 1190 1308 1606 1311
rect 1610 1308 1729 1311
rect 1738 1308 1774 1311
rect 1866 1308 1878 1311
rect 1898 1308 1934 1311
rect 2098 1308 2118 1311
rect 2122 1308 2134 1311
rect 2202 1308 2318 1311
rect 2354 1308 2366 1311
rect 2378 1308 2454 1311
rect 2474 1308 2478 1311
rect 2586 1308 2606 1311
rect 2674 1308 2782 1311
rect 2790 1308 2990 1311
rect 3090 1308 3190 1311
rect 3362 1308 3446 1311
rect 14 1302 17 1308
rect 992 1303 994 1307
rect 998 1303 1001 1307
rect 1006 1303 1008 1307
rect 322 1298 374 1301
rect 394 1298 406 1301
rect 666 1298 702 1301
rect 714 1298 734 1301
rect 754 1298 846 1301
rect 874 1298 926 1301
rect 930 1298 974 1301
rect 1018 1298 1078 1301
rect 1130 1298 1142 1301
rect 1194 1298 1334 1301
rect 1386 1298 1390 1301
rect 1426 1298 1582 1301
rect 1594 1298 1710 1301
rect 1726 1301 1729 1308
rect 1726 1298 1750 1301
rect 1758 1298 1774 1301
rect 1782 1301 1785 1308
rect 1886 1302 1889 1308
rect 2024 1303 2026 1307
rect 2030 1303 2033 1307
rect 2038 1303 2040 1307
rect 1782 1298 1854 1301
rect 1906 1298 1910 1301
rect 1954 1298 1974 1301
rect 1978 1298 2014 1301
rect 2090 1298 2126 1301
rect 2186 1298 2206 1301
rect 2210 1298 2222 1301
rect 2266 1298 2302 1301
rect 2318 1301 2321 1308
rect 2318 1298 2390 1301
rect 2434 1298 2606 1301
rect 2790 1301 2793 1308
rect 3040 1303 3042 1307
rect 3046 1303 3049 1307
rect 3054 1303 3056 1307
rect 2610 1298 2793 1301
rect 2834 1298 2838 1301
rect 2850 1298 2854 1301
rect 2882 1298 3014 1301
rect 3018 1298 3030 1301
rect 3090 1298 3254 1301
rect 3258 1298 3366 1301
rect 3378 1298 3462 1301
rect 14 1288 70 1291
rect 346 1288 454 1291
rect 490 1288 1030 1291
rect 1042 1288 1054 1291
rect 1094 1288 1158 1291
rect 1194 1288 1206 1291
rect 1270 1288 1278 1291
rect 1298 1288 1302 1291
rect 1326 1288 1334 1291
rect 1338 1288 1366 1291
rect 1378 1288 1398 1291
rect 1514 1288 1542 1291
rect 1562 1288 1566 1291
rect 1578 1288 1582 1291
rect 1594 1288 1598 1291
rect 1618 1288 1718 1291
rect 1758 1291 1761 1298
rect 1722 1288 1761 1291
rect 1770 1288 1798 1291
rect 1810 1288 1910 1291
rect 1930 1288 1950 1291
rect 1978 1288 2110 1291
rect 2146 1288 2174 1291
rect 2194 1288 2206 1291
rect 2218 1288 2246 1291
rect 2298 1288 2382 1291
rect 2442 1288 2454 1291
rect 2458 1288 2462 1291
rect 2510 1288 2518 1291
rect 2522 1288 2590 1291
rect 2618 1288 3142 1291
rect 3146 1288 3254 1291
rect 3274 1288 3318 1291
rect 3418 1288 3478 1291
rect 14 1282 17 1288
rect 166 1282 169 1288
rect 1094 1282 1097 1288
rect 1254 1282 1257 1288
rect 1262 1282 1265 1288
rect 2286 1282 2289 1288
rect 2406 1282 2409 1288
rect 138 1278 142 1281
rect 170 1278 198 1281
rect 258 1278 278 1281
rect 338 1278 350 1281
rect 362 1278 398 1281
rect 426 1278 430 1281
rect 446 1278 617 1281
rect 170 1268 190 1271
rect 194 1268 209 1271
rect 218 1268 294 1271
rect 298 1268 318 1271
rect 370 1268 382 1271
rect 402 1268 414 1271
rect 438 1271 441 1278
rect 418 1268 441 1271
rect 446 1272 449 1278
rect 614 1272 617 1278
rect 634 1278 790 1281
rect 810 1278 854 1281
rect 898 1278 926 1281
rect 938 1278 966 1281
rect 978 1278 1070 1281
rect 1170 1278 1222 1281
rect 1282 1278 1774 1281
rect 1826 1278 1830 1281
rect 1850 1278 1862 1281
rect 1874 1278 1966 1281
rect 2018 1278 2030 1281
rect 2082 1278 2118 1281
rect 2126 1278 2262 1281
rect 2322 1278 2382 1281
rect 2386 1278 2390 1281
rect 2418 1278 2470 1281
rect 2530 1278 2534 1281
rect 2762 1278 2918 1281
rect 2922 1278 2926 1281
rect 2986 1278 3001 1281
rect 3194 1278 3214 1281
rect 3254 1281 3257 1288
rect 3254 1278 3374 1281
rect 3410 1278 3414 1281
rect 622 1272 625 1278
rect 630 1272 633 1278
rect 1838 1272 1841 1278
rect 498 1268 566 1271
rect 586 1268 598 1271
rect 658 1268 718 1271
rect 746 1268 750 1271
rect 802 1268 822 1271
rect 842 1268 846 1271
rect 970 1268 974 1271
rect 986 1268 1006 1271
rect 1018 1268 1038 1271
rect 1082 1268 1094 1271
rect 1106 1268 1126 1271
rect 1162 1268 1185 1271
rect 1226 1268 1246 1271
rect 1250 1268 1286 1271
rect 1314 1268 1334 1271
rect 1338 1268 1342 1271
rect 1362 1268 1422 1271
rect 1434 1268 1438 1271
rect 1466 1268 1550 1271
rect 1630 1268 1638 1271
rect 1650 1268 1662 1271
rect 1674 1268 1678 1271
rect 1706 1268 1710 1271
rect 1802 1268 1838 1271
rect 1850 1268 1894 1271
rect 1906 1268 1910 1271
rect 1938 1268 1942 1271
rect 1954 1268 1982 1271
rect 2002 1268 2022 1271
rect 2034 1268 2086 1271
rect 2126 1271 2129 1278
rect 2122 1268 2129 1271
rect 2138 1268 2142 1271
rect 2162 1268 2166 1271
rect 2210 1268 2238 1271
rect 2250 1268 2374 1271
rect 2394 1268 2494 1271
rect 2626 1268 2630 1271
rect 2642 1268 2646 1271
rect 2706 1268 2782 1271
rect 2786 1268 2846 1271
rect 2850 1268 2862 1271
rect 2882 1268 2894 1271
rect 2898 1268 2934 1271
rect 2966 1271 2969 1278
rect 2998 1272 3001 1278
rect 2966 1268 2974 1271
rect 3010 1268 3038 1271
rect 3042 1268 3110 1271
rect 3114 1268 3150 1271
rect 3170 1268 3342 1271
rect 3426 1268 3446 1271
rect 3450 1268 3486 1271
rect 3490 1268 3558 1271
rect 18 1258 62 1261
rect 90 1258 102 1261
rect 182 1258 190 1261
rect 194 1258 198 1261
rect 206 1261 209 1268
rect 350 1261 353 1268
rect 206 1258 430 1261
rect 438 1261 441 1268
rect 438 1258 558 1261
rect 606 1261 609 1268
rect 782 1262 785 1268
rect 870 1262 873 1268
rect 1062 1262 1065 1268
rect 1070 1262 1073 1268
rect 1102 1262 1105 1268
rect 594 1258 609 1261
rect 618 1258 638 1261
rect 650 1258 726 1261
rect 802 1258 806 1261
rect 818 1258 838 1261
rect 842 1258 854 1261
rect 922 1258 942 1261
rect 954 1258 982 1261
rect 1026 1258 1030 1261
rect 1162 1258 1174 1261
rect 1182 1261 1185 1268
rect 1182 1258 1206 1261
rect 1218 1258 1286 1261
rect 1302 1258 1318 1261
rect 1346 1258 1353 1261
rect 1378 1258 1446 1261
rect 1482 1258 1550 1261
rect 1562 1258 1566 1261
rect 1578 1258 1598 1261
rect 1610 1258 1622 1261
rect 1630 1261 1633 1268
rect 1734 1262 1737 1268
rect 1758 1262 1761 1268
rect 1626 1258 1633 1261
rect 1642 1258 1649 1261
rect 1674 1258 1686 1261
rect 1706 1258 1710 1261
rect 1746 1258 1750 1261
rect 1826 1258 1870 1261
rect 1882 1258 1894 1261
rect 1906 1258 1910 1261
rect 2094 1261 2097 1268
rect 1946 1258 2097 1261
rect 2114 1258 2158 1261
rect 2222 1258 2270 1261
rect 2290 1258 2422 1261
rect 2442 1258 2446 1261
rect 2450 1258 2462 1261
rect 2498 1258 2590 1261
rect 2690 1258 2718 1261
rect 2746 1258 2814 1261
rect 2858 1258 2902 1261
rect 2922 1258 2926 1261
rect 2978 1258 3014 1261
rect 3018 1258 3054 1261
rect 3122 1258 3182 1261
rect 3250 1258 3278 1261
rect 3282 1258 3310 1261
rect 3346 1258 3358 1261
rect 3402 1258 3417 1261
rect 3426 1258 3430 1261
rect 718 1252 721 1258
rect 34 1248 134 1251
rect 194 1248 198 1251
rect 226 1248 230 1251
rect 242 1248 246 1251
rect 290 1248 294 1251
rect 314 1248 374 1251
rect 402 1248 406 1251
rect 478 1248 486 1251
rect 490 1248 654 1251
rect 690 1248 694 1251
rect 770 1248 1086 1251
rect 1094 1251 1097 1258
rect 1094 1248 1126 1251
rect 1146 1248 1166 1251
rect 1226 1248 1238 1251
rect 1302 1251 1305 1258
rect 1350 1252 1353 1258
rect 1646 1252 1649 1258
rect 1282 1248 1305 1251
rect 1314 1248 1318 1251
rect 1330 1248 1342 1251
rect 1370 1248 1414 1251
rect 1426 1248 1486 1251
rect 1546 1248 1574 1251
rect 1586 1248 1638 1251
rect 1654 1248 1806 1251
rect 1826 1248 1846 1251
rect 1858 1248 2166 1251
rect 2222 1251 2225 1258
rect 2186 1248 2225 1251
rect 2234 1248 2326 1251
rect 2346 1248 2350 1251
rect 2478 1251 2481 1258
rect 2718 1252 2721 1258
rect 2478 1248 2550 1251
rect 2578 1248 2614 1251
rect 2634 1248 2638 1251
rect 2658 1248 2710 1251
rect 2770 1248 2774 1251
rect 2834 1248 2838 1251
rect 2942 1251 2945 1258
rect 2890 1248 2945 1251
rect 2962 1248 3134 1251
rect 3194 1248 3198 1251
rect 3282 1248 3286 1251
rect 3290 1248 3350 1251
rect 3378 1248 3390 1251
rect 3414 1251 3417 1258
rect 3414 1248 3494 1251
rect 3590 1248 3594 1252
rect 374 1242 377 1248
rect 202 1238 214 1241
rect 218 1238 238 1241
rect 322 1238 334 1241
rect 422 1241 425 1248
rect 422 1238 438 1241
rect 458 1238 902 1241
rect 930 1238 982 1241
rect 1026 1238 1078 1241
rect 1130 1238 1214 1241
rect 1246 1241 1249 1248
rect 1246 1238 1278 1241
rect 1298 1238 1318 1241
rect 1338 1238 1606 1241
rect 1654 1241 1657 1248
rect 1618 1238 1657 1241
rect 1674 1238 1766 1241
rect 1850 1238 1990 1241
rect 1998 1238 2022 1241
rect 2058 1238 2062 1241
rect 2082 1238 2094 1241
rect 2106 1238 2150 1241
rect 2162 1238 2198 1241
rect 2274 1238 2414 1241
rect 2434 1238 2486 1241
rect 2562 1238 2726 1241
rect 2746 1238 2750 1241
rect 2778 1238 2926 1241
rect 2970 1238 3070 1241
rect 3590 1241 3593 1248
rect 3154 1238 3593 1241
rect 74 1228 614 1231
rect 642 1228 646 1231
rect 778 1228 798 1231
rect 858 1228 1038 1231
rect 1058 1228 1094 1231
rect 1102 1228 1190 1231
rect 1210 1228 1222 1231
rect 1266 1228 1390 1231
rect 1394 1228 1414 1231
rect 1426 1228 1454 1231
rect 1474 1228 1478 1231
rect 1482 1228 1550 1231
rect 1562 1228 1654 1231
rect 1666 1228 1694 1231
rect 1742 1228 1750 1231
rect 1754 1228 1774 1231
rect 1814 1231 1817 1238
rect 1794 1228 1817 1231
rect 1834 1228 1985 1231
rect 1998 1231 2001 1238
rect 1994 1228 2001 1231
rect 2030 1228 2134 1231
rect 2146 1228 2150 1231
rect 2194 1228 2198 1231
rect 2206 1231 2209 1238
rect 2206 1228 2286 1231
rect 2298 1228 2302 1231
rect 2330 1228 2598 1231
rect 2610 1228 2806 1231
rect 2810 1228 2814 1231
rect 2926 1231 2929 1238
rect 2926 1228 3126 1231
rect 3326 1228 3342 1231
rect 146 1218 518 1221
rect 570 1218 646 1221
rect 686 1221 689 1228
rect 686 1218 862 1221
rect 1102 1221 1105 1228
rect 1198 1222 1201 1228
rect 906 1218 1105 1221
rect 1114 1218 1166 1221
rect 1206 1218 1214 1221
rect 1218 1218 1286 1221
rect 1298 1218 1302 1221
rect 1314 1218 1326 1221
rect 1338 1218 1342 1221
rect 1362 1218 1414 1221
rect 1426 1218 1881 1221
rect 1890 1218 1894 1221
rect 1922 1218 1966 1221
rect 1982 1221 1985 1228
rect 2030 1221 2033 1228
rect 3326 1222 3329 1228
rect 1970 1218 1977 1221
rect 1982 1218 2033 1221
rect 2042 1218 2046 1221
rect 2058 1218 2230 1221
rect 2274 1218 2302 1221
rect 2330 1218 2422 1221
rect 2434 1218 2494 1221
rect 2570 1218 2798 1221
rect 2922 1218 3294 1221
rect 82 1208 310 1211
rect 322 1208 470 1211
rect 518 1211 521 1218
rect 518 1208 582 1211
rect 786 1208 1025 1211
rect 1042 1208 1390 1211
rect 1434 1208 1470 1211
rect 1482 1208 1494 1211
rect 1562 1208 1630 1211
rect 1642 1208 1830 1211
rect 1842 1208 1870 1211
rect 1878 1211 1881 1218
rect 1878 1208 1910 1211
rect 1914 1208 2014 1211
rect 2026 1208 2046 1211
rect 2082 1208 2118 1211
rect 2138 1208 2334 1211
rect 2354 1208 2446 1211
rect 2634 1208 3022 1211
rect 3074 1208 3126 1211
rect 480 1203 482 1207
rect 486 1203 489 1207
rect 494 1203 496 1207
rect 1022 1202 1025 1208
rect 1512 1203 1514 1207
rect 1518 1203 1521 1207
rect 1526 1203 1528 1207
rect 2536 1203 2538 1207
rect 2542 1203 2545 1207
rect 2550 1203 2552 1207
rect 266 1198 462 1201
rect 506 1198 726 1201
rect 746 1198 750 1201
rect 874 1198 934 1201
rect 954 1198 958 1201
rect 1002 1198 1009 1201
rect 1042 1198 1054 1201
rect 1066 1198 1070 1201
rect 1082 1198 1198 1201
rect 1242 1198 1254 1201
rect 1306 1198 1310 1201
rect 1322 1198 1334 1201
rect 1394 1198 1462 1201
rect 1558 1198 1838 1201
rect 1846 1198 1998 1201
rect 2002 1198 2014 1201
rect 2018 1198 2070 1201
rect 2074 1198 2134 1201
rect 2138 1198 2206 1201
rect 2218 1198 2526 1201
rect 2634 1198 2638 1201
rect 2946 1198 2966 1201
rect 3018 1198 3182 1201
rect 3186 1198 3254 1201
rect 990 1192 993 1198
rect 138 1188 206 1191
rect 238 1188 390 1191
rect 450 1188 542 1191
rect 554 1188 630 1191
rect 634 1188 665 1191
rect 778 1188 814 1191
rect 938 1188 942 1191
rect 954 1188 966 1191
rect 1006 1191 1009 1198
rect 1006 1188 1110 1191
rect 1130 1188 1182 1191
rect 1186 1188 1262 1191
rect 1322 1188 1326 1191
rect 1410 1188 1446 1191
rect 1558 1191 1561 1198
rect 1846 1192 1849 1198
rect 1498 1188 1561 1191
rect 1570 1188 1598 1191
rect 1634 1188 1646 1191
rect 1658 1188 1670 1191
rect 1714 1188 1798 1191
rect 1802 1188 1846 1191
rect 1858 1188 1942 1191
rect 1962 1188 2030 1191
rect 2050 1188 2118 1191
rect 2126 1188 2238 1191
rect 2242 1188 2414 1191
rect 2642 1188 2710 1191
rect 3066 1188 3158 1191
rect 238 1182 241 1188
rect 274 1178 318 1181
rect 398 1181 401 1188
rect 322 1178 401 1181
rect 530 1178 654 1181
rect 662 1181 665 1188
rect 662 1178 1102 1181
rect 1178 1178 1214 1181
rect 1242 1178 1334 1181
rect 1350 1181 1353 1188
rect 2126 1182 2129 1188
rect 1350 1178 1390 1181
rect 1418 1178 1454 1181
rect 1466 1178 1750 1181
rect 1762 1178 1870 1181
rect 1882 1178 1918 1181
rect 1930 1178 1998 1181
rect 2066 1178 2086 1181
rect 2146 1178 2374 1181
rect 2386 1178 2430 1181
rect 2450 1178 2582 1181
rect 2642 1178 2646 1181
rect 2870 1181 2873 1188
rect 2786 1178 2873 1181
rect 66 1168 94 1171
rect 210 1168 222 1171
rect 290 1168 942 1171
rect 1158 1171 1161 1178
rect 1130 1168 1161 1171
rect 1210 1168 1238 1171
rect 1274 1168 1366 1171
rect 1370 1168 1430 1171
rect 1434 1168 1462 1171
rect 1474 1168 1478 1171
rect 1490 1168 1494 1171
rect 1538 1168 1582 1171
rect 1602 1168 1713 1171
rect 1722 1168 1886 1171
rect 1902 1168 1910 1171
rect 1914 1168 1918 1171
rect 1930 1168 2158 1171
rect 2170 1168 2198 1171
rect 2202 1168 2334 1171
rect 2506 1168 2574 1171
rect 2586 1168 2614 1171
rect 2618 1168 2622 1171
rect 2722 1168 2750 1171
rect 2762 1168 2790 1171
rect 2962 1168 3086 1171
rect 3098 1168 3174 1171
rect 3178 1168 3302 1171
rect 3306 1168 3310 1171
rect 3398 1171 3401 1178
rect 3398 1168 3446 1171
rect 3590 1171 3594 1172
rect 3562 1168 3594 1171
rect 166 1162 169 1168
rect 1246 1162 1249 1168
rect 98 1158 102 1161
rect 290 1158 510 1161
rect 562 1158 606 1161
rect 738 1158 766 1161
rect 802 1158 822 1161
rect 890 1158 1158 1161
rect 1266 1158 1286 1161
rect 1322 1158 1462 1161
rect 1514 1158 1622 1161
rect 1650 1158 1654 1161
rect 1674 1158 1686 1161
rect 1710 1161 1713 1168
rect 1710 1158 1718 1161
rect 1722 1158 1750 1161
rect 1778 1158 1782 1161
rect 1810 1158 1814 1161
rect 1826 1158 1833 1161
rect 1866 1158 1958 1161
rect 1970 1158 1982 1161
rect 2002 1158 2054 1161
rect 2066 1158 2174 1161
rect 2242 1158 2310 1161
rect 2322 1158 2406 1161
rect 2418 1158 2678 1161
rect 2682 1158 2782 1161
rect 2818 1158 2982 1161
rect 3026 1158 3030 1161
rect 3378 1158 3406 1161
rect 3422 1158 3462 1161
rect 678 1152 681 1158
rect 34 1148 102 1151
rect 202 1148 270 1151
rect 322 1148 342 1151
rect 418 1148 438 1151
rect 522 1148 534 1151
rect 610 1148 649 1151
rect 698 1148 702 1151
rect 722 1148 726 1151
rect 738 1148 750 1151
rect 810 1148 822 1151
rect 826 1148 830 1151
rect 838 1151 841 1158
rect 846 1151 849 1158
rect 838 1148 849 1151
rect 970 1148 998 1151
rect 1018 1148 1022 1151
rect 1090 1148 1142 1151
rect 1174 1151 1177 1158
rect 1830 1152 1833 1158
rect 1174 1148 1182 1151
rect 1226 1148 1230 1151
rect 1234 1148 1246 1151
rect 1250 1148 1286 1151
rect 1314 1148 1478 1151
rect 1506 1148 1510 1151
rect 1530 1148 1534 1151
rect 1570 1148 1593 1151
rect 398 1142 401 1148
rect 646 1142 649 1148
rect 750 1142 753 1148
rect 1054 1142 1057 1148
rect 1294 1142 1297 1148
rect 1302 1142 1305 1148
rect 1590 1142 1593 1148
rect 1634 1148 1646 1151
rect 1650 1148 1686 1151
rect 1698 1148 1718 1151
rect 1722 1148 1726 1151
rect 1746 1148 1758 1151
rect 1778 1148 1806 1151
rect 1866 1148 1870 1151
rect 1890 1148 1982 1151
rect 1990 1151 1993 1158
rect 1990 1148 1998 1151
rect 2026 1148 2054 1151
rect 2058 1148 2142 1151
rect 2218 1148 2230 1151
rect 2238 1148 2254 1151
rect 2266 1148 2270 1151
rect 2370 1148 2382 1151
rect 2510 1148 2614 1151
rect 2706 1148 2806 1151
rect 2810 1148 2862 1151
rect 3114 1148 3150 1151
rect 3178 1148 3182 1151
rect 3194 1148 3342 1151
rect 3366 1151 3369 1158
rect 3422 1151 3425 1158
rect 3366 1148 3425 1151
rect 3434 1148 3526 1151
rect 3590 1151 3594 1152
rect 3562 1148 3594 1151
rect 1606 1142 1609 1148
rect 2174 1142 2177 1148
rect 50 1138 73 1141
rect 98 1138 113 1141
rect 6 1132 9 1138
rect 70 1132 73 1138
rect 110 1132 113 1138
rect 146 1138 182 1141
rect 186 1138 206 1141
rect 426 1138 526 1141
rect 658 1138 694 1141
rect 762 1138 798 1141
rect 818 1138 838 1141
rect 850 1138 854 1141
rect 866 1138 878 1141
rect 882 1138 910 1141
rect 922 1138 934 1141
rect 938 1138 966 1141
rect 1026 1138 1038 1141
rect 1082 1138 1182 1141
rect 1210 1138 1230 1141
rect 1342 1138 1350 1141
rect 1354 1138 1366 1141
rect 1370 1138 1414 1141
rect 1418 1138 1438 1141
rect 1442 1138 1486 1141
rect 1562 1138 1582 1141
rect 1634 1138 1638 1141
rect 1658 1138 1702 1141
rect 1730 1138 1734 1141
rect 1754 1138 1774 1141
rect 1802 1138 1854 1141
rect 1870 1138 1977 1141
rect 1986 1138 1990 1141
rect 2026 1138 2070 1141
rect 2082 1138 2102 1141
rect 2122 1138 2142 1141
rect 2198 1141 2201 1148
rect 2238 1141 2241 1148
rect 2510 1142 2513 1148
rect 2198 1138 2241 1141
rect 2258 1138 2398 1141
rect 2402 1138 2478 1141
rect 2522 1138 2526 1141
rect 2578 1138 2662 1141
rect 2682 1138 2694 1141
rect 2706 1138 2710 1141
rect 2738 1138 2742 1141
rect 2754 1138 2846 1141
rect 2882 1138 2886 1141
rect 2890 1138 2934 1141
rect 2962 1138 2966 1141
rect 3002 1138 3094 1141
rect 3114 1138 3134 1141
rect 3154 1138 3214 1141
rect 3306 1138 3326 1141
rect 3346 1138 3374 1141
rect 134 1132 137 1138
rect 742 1132 745 1138
rect 1238 1132 1241 1138
rect 410 1128 462 1131
rect 674 1128 686 1131
rect 754 1128 774 1131
rect 782 1128 790 1131
rect 794 1128 886 1131
rect 946 1128 950 1131
rect 1034 1128 1062 1131
rect 1170 1128 1190 1131
rect 1194 1128 1238 1131
rect 1282 1128 1302 1131
rect 1342 1131 1345 1138
rect 1550 1132 1553 1138
rect 1614 1132 1617 1138
rect 1338 1128 1345 1131
rect 1354 1128 1358 1131
rect 1370 1128 1422 1131
rect 1434 1128 1478 1131
rect 1578 1128 1606 1131
rect 1642 1128 1646 1131
rect 1666 1128 1702 1131
rect 1754 1128 1782 1131
rect 1794 1128 1798 1131
rect 1870 1131 1873 1138
rect 1834 1128 1873 1131
rect 1882 1128 1926 1131
rect 1938 1128 1942 1131
rect 1974 1131 1977 1138
rect 1974 1128 1998 1131
rect 2006 1131 2009 1138
rect 3382 1132 3385 1138
rect 2006 1128 2206 1131
rect 2210 1128 2238 1131
rect 2314 1128 2454 1131
rect 2482 1128 2486 1131
rect 2522 1128 2526 1131
rect 2546 1128 2550 1131
rect 2722 1128 2758 1131
rect 2778 1128 2822 1131
rect 2826 1128 2862 1131
rect 2870 1128 2902 1131
rect 2906 1128 2950 1131
rect 3002 1128 3014 1131
rect 3034 1128 3110 1131
rect 3186 1128 3198 1131
rect 3218 1128 3230 1131
rect 3242 1128 3358 1131
rect 910 1122 913 1128
rect 926 1122 929 1128
rect 1326 1122 1329 1128
rect 2662 1122 2665 1128
rect 10 1118 254 1121
rect 274 1118 438 1121
rect 570 1118 766 1121
rect 778 1118 830 1121
rect 834 1118 862 1121
rect 946 1118 974 1121
rect 986 1118 1118 1121
rect 1186 1118 1262 1121
rect 1278 1118 1318 1121
rect 1346 1118 1606 1121
rect 1626 1118 1662 1121
rect 1706 1118 1814 1121
rect 1834 1118 1862 1121
rect 1890 1118 1910 1121
rect 1938 1118 2006 1121
rect 2014 1118 2038 1121
rect 2074 1118 2318 1121
rect 2370 1118 2406 1121
rect 2870 1121 2873 1128
rect 2698 1118 2873 1121
rect 2882 1118 3166 1121
rect 3242 1118 3262 1121
rect 3306 1118 3326 1121
rect 178 1108 454 1111
rect 506 1108 726 1111
rect 738 1108 822 1111
rect 858 1108 950 1111
rect 1026 1108 1110 1111
rect 1122 1108 1206 1111
rect 1218 1108 1222 1111
rect 1278 1111 1281 1118
rect 1258 1108 1281 1111
rect 1290 1108 1926 1111
rect 1962 1108 1982 1111
rect 2014 1111 2017 1118
rect 3278 1112 3281 1118
rect 1994 1108 2017 1111
rect 2074 1108 2102 1111
rect 2114 1108 2126 1111
rect 2138 1108 2486 1111
rect 2490 1108 2774 1111
rect 2802 1108 2830 1111
rect 2898 1108 2998 1111
rect 3162 1108 3214 1111
rect 992 1103 994 1107
rect 998 1103 1001 1107
rect 1006 1103 1008 1107
rect 2024 1103 2026 1107
rect 2030 1103 2033 1107
rect 2038 1103 2040 1107
rect 3040 1103 3042 1107
rect 3046 1103 3049 1107
rect 3054 1103 3056 1107
rect 3310 1102 3313 1108
rect 3494 1102 3497 1108
rect 74 1098 118 1101
rect 378 1098 390 1101
rect 434 1098 518 1101
rect 522 1098 534 1101
rect 594 1098 622 1101
rect 642 1098 654 1101
rect 698 1098 870 1101
rect 914 1098 926 1101
rect 930 1098 958 1101
rect 1058 1098 1078 1101
rect 1178 1098 1241 1101
rect 1290 1098 1294 1101
rect 1306 1098 1366 1101
rect 1402 1098 1406 1101
rect 1442 1098 1446 1101
rect 1474 1098 1486 1101
rect 1554 1098 1638 1101
rect 1666 1098 1710 1101
rect 1722 1098 1726 1101
rect 1778 1098 1798 1101
rect 1810 1098 1814 1101
rect 1962 1098 1998 1101
rect 2050 1098 2222 1101
rect 2250 1098 2262 1101
rect 2314 1098 2350 1101
rect 2530 1098 2558 1101
rect 2562 1098 2718 1101
rect 2738 1098 2774 1101
rect 2810 1098 2814 1101
rect 2906 1098 3006 1101
rect 3010 1098 3030 1101
rect 3066 1098 3126 1101
rect 3130 1098 3214 1101
rect 398 1088 406 1091
rect 410 1088 478 1091
rect 482 1088 558 1091
rect 586 1088 774 1091
rect 826 1088 878 1091
rect 898 1088 942 1091
rect 954 1088 990 1091
rect 1002 1088 1014 1091
rect 1034 1088 1086 1091
rect 1122 1088 1142 1091
rect 1146 1088 1150 1091
rect 1194 1088 1230 1091
rect 1238 1091 1241 1098
rect 1894 1092 1897 1098
rect 1238 1088 1270 1091
rect 1282 1088 1310 1091
rect 1322 1088 1374 1091
rect 1378 1088 1526 1091
rect 1538 1088 1542 1091
rect 1554 1088 1582 1091
rect 1594 1088 1654 1091
rect 1706 1088 1830 1091
rect 1866 1088 1886 1091
rect 2006 1088 2014 1091
rect 2018 1088 2046 1091
rect 2066 1088 2086 1091
rect 2122 1088 2150 1091
rect 2186 1088 2246 1091
rect 2266 1088 2294 1091
rect 2354 1088 2366 1091
rect 2402 1088 2430 1091
rect 2498 1088 2510 1091
rect 2514 1088 2998 1091
rect 3034 1088 3086 1091
rect 3282 1088 3286 1091
rect 3294 1091 3297 1098
rect 3294 1088 3382 1091
rect 3434 1088 3518 1091
rect 86 1082 89 1088
rect 42 1078 78 1081
rect 346 1078 462 1081
rect 626 1078 662 1081
rect 690 1078 886 1081
rect 970 1078 1110 1081
rect 1130 1078 1446 1081
rect 1466 1078 1630 1081
rect 1658 1078 1670 1081
rect 1686 1081 1689 1088
rect 1838 1082 1841 1088
rect 2062 1082 2065 1088
rect 1686 1078 1726 1081
rect 1738 1078 1766 1081
rect 1770 1078 1774 1081
rect 1810 1078 1830 1081
rect 1850 1078 1878 1081
rect 1890 1078 1910 1081
rect 1938 1078 1966 1081
rect 1978 1078 2046 1081
rect 2074 1078 2182 1081
rect 2186 1078 2206 1081
rect 2218 1078 2230 1081
rect 2306 1078 2310 1081
rect 2370 1078 2382 1081
rect 2406 1078 2558 1081
rect 2618 1078 2622 1081
rect 2658 1078 2686 1081
rect 2706 1078 2718 1081
rect 2722 1078 2726 1081
rect 2842 1078 2846 1081
rect 3122 1078 3150 1081
rect 3162 1078 3206 1081
rect 3226 1078 3334 1081
rect 3590 1078 3594 1082
rect 66 1068 134 1071
rect 154 1068 182 1071
rect 186 1068 190 1071
rect 298 1068 350 1071
rect 362 1068 366 1071
rect 410 1068 422 1071
rect 474 1068 513 1071
rect 570 1068 590 1071
rect 610 1068 622 1071
rect 674 1068 718 1071
rect 722 1068 742 1071
rect 746 1068 758 1071
rect 786 1068 798 1071
rect 810 1068 830 1071
rect 850 1068 966 1071
rect 978 1068 982 1071
rect 1090 1068 1110 1071
rect 1138 1068 1246 1071
rect 1250 1068 1254 1071
rect 1266 1068 1318 1071
rect 1338 1068 1374 1071
rect 1386 1068 1430 1071
rect 1538 1068 1542 1071
rect 1578 1068 1590 1071
rect 1610 1068 1622 1071
rect 1654 1071 1657 1078
rect 1634 1068 1649 1071
rect 1654 1068 1662 1071
rect 1682 1068 1694 1071
rect 1714 1068 1718 1071
rect 1750 1068 1766 1071
rect 1794 1068 1878 1071
rect 1882 1068 1902 1071
rect 1906 1068 1950 1071
rect 1978 1068 1982 1071
rect 1994 1068 2006 1071
rect 2010 1068 2038 1071
rect 2050 1068 2086 1071
rect 2098 1068 2110 1071
rect 2122 1068 2190 1071
rect 2218 1068 2230 1071
rect 2406 1071 2409 1078
rect 2910 1072 2913 1078
rect 2926 1072 2929 1078
rect 2266 1068 2409 1071
rect 2430 1068 2438 1071
rect 2546 1068 2550 1071
rect 2618 1068 2665 1071
rect 2690 1068 2718 1071
rect 2810 1068 2894 1071
rect 2938 1068 2942 1071
rect 3002 1068 3166 1071
rect 3186 1068 3246 1071
rect 3590 1071 3593 1078
rect 3250 1068 3593 1071
rect 510 1062 513 1068
rect 1022 1062 1025 1068
rect 1126 1062 1129 1068
rect 18 1058 118 1061
rect 122 1058 142 1061
rect 178 1058 222 1061
rect 242 1058 294 1061
rect 298 1058 334 1061
rect 354 1058 390 1061
rect 394 1058 422 1061
rect 426 1058 438 1061
rect 458 1058 470 1061
rect 514 1058 518 1061
rect 554 1058 582 1061
rect 586 1058 606 1061
rect 626 1058 638 1061
rect 658 1058 694 1061
rect 714 1058 718 1061
rect 754 1058 782 1061
rect 794 1058 830 1061
rect 842 1058 950 1061
rect 994 1058 1006 1061
rect 1034 1058 1038 1061
rect 1050 1058 1054 1061
rect 1066 1058 1070 1061
rect 1106 1058 1110 1061
rect 1178 1058 1190 1061
rect 1194 1058 1206 1061
rect 1218 1058 1222 1061
rect 1234 1058 1446 1061
rect 1506 1058 1510 1061
rect 1530 1058 1606 1061
rect 1646 1061 1649 1068
rect 1750 1061 1753 1068
rect 2414 1062 2417 1068
rect 2430 1062 2433 1068
rect 2662 1062 2665 1068
rect 1646 1058 1753 1061
rect 1762 1058 1894 1061
rect 1906 1058 1998 1061
rect 2090 1058 2094 1061
rect 2162 1058 2166 1061
rect 2290 1058 2318 1061
rect 2338 1058 2374 1061
rect 2690 1058 2710 1061
rect 2734 1058 2766 1061
rect 2786 1058 2878 1061
rect 2946 1058 2958 1061
rect 2994 1058 3062 1061
rect 3106 1058 3126 1061
rect 3174 1061 3177 1068
rect 3174 1058 3230 1061
rect 3290 1058 3326 1061
rect 3330 1058 3361 1061
rect 3386 1058 3406 1061
rect 1630 1052 1633 1058
rect 2326 1052 2329 1058
rect 2710 1052 2713 1058
rect 2734 1052 2737 1058
rect 18 1048 22 1051
rect 74 1048 78 1051
rect 114 1048 150 1051
rect 154 1048 662 1051
rect 682 1048 806 1051
rect 818 1048 822 1051
rect 858 1048 862 1051
rect 866 1048 878 1051
rect 890 1048 918 1051
rect 930 1048 942 1051
rect 994 1048 1038 1051
rect 1058 1048 1070 1051
rect 1162 1048 1206 1051
rect 1242 1048 1254 1051
rect 1266 1048 1278 1051
rect 1322 1048 1398 1051
rect 1410 1048 1510 1051
rect 1594 1048 1614 1051
rect 1650 1048 1654 1051
rect 1666 1048 1670 1051
rect 1706 1048 1742 1051
rect 1746 1048 1758 1051
rect 1770 1048 1886 1051
rect 1906 1048 1918 1051
rect 1926 1048 1942 1051
rect 1970 1048 1993 1051
rect 2002 1048 2062 1051
rect 2082 1048 2086 1051
rect 2098 1048 2110 1051
rect 2258 1048 2278 1051
rect 2290 1048 2294 1051
rect 2306 1048 2310 1051
rect 2402 1048 2558 1051
rect 2850 1048 2854 1051
rect 2874 1048 2902 1051
rect 2918 1051 2921 1058
rect 3358 1052 3361 1058
rect 2918 1048 2942 1051
rect 3066 1048 3150 1051
rect 3154 1048 3198 1051
rect 3202 1048 3254 1051
rect 3338 1048 3350 1051
rect 3370 1048 3374 1051
rect 3402 1048 3462 1051
rect 3590 1051 3594 1052
rect 3562 1048 3594 1051
rect 1694 1042 1697 1048
rect 10 1038 30 1041
rect 98 1038 118 1041
rect 126 1038 174 1041
rect 234 1038 278 1041
rect 354 1038 438 1041
rect 450 1038 502 1041
rect 514 1038 526 1041
rect 578 1038 582 1041
rect 594 1038 606 1041
rect 658 1038 662 1041
rect 730 1038 1110 1041
rect 1178 1038 1286 1041
rect 1290 1038 1294 1041
rect 1330 1038 1342 1041
rect 1354 1038 1358 1041
rect 1530 1038 1686 1041
rect 1714 1038 1878 1041
rect 1926 1041 1929 1048
rect 1906 1038 1929 1041
rect 1946 1038 1966 1041
rect 1990 1041 1993 1048
rect 1990 1038 2166 1041
rect 2174 1041 2177 1048
rect 2174 1038 2222 1041
rect 2234 1038 2302 1041
rect 2314 1038 2494 1041
rect 2594 1038 2742 1041
rect 2746 1038 2782 1041
rect 2802 1038 3086 1041
rect 3090 1038 3182 1041
rect 3186 1038 3198 1041
rect 3218 1038 3318 1041
rect 3322 1038 3350 1041
rect 3410 1038 3430 1041
rect 126 1032 129 1038
rect 206 1032 209 1038
rect 378 1028 590 1031
rect 778 1028 886 1031
rect 938 1028 950 1031
rect 1098 1028 1198 1031
rect 1258 1028 1406 1031
rect 1426 1028 1430 1031
rect 1466 1028 1558 1031
rect 1570 1028 1814 1031
rect 1882 1028 2150 1031
rect 2154 1028 2446 1031
rect 2522 1028 2806 1031
rect 2818 1028 2918 1031
rect 2946 1028 3022 1031
rect 3050 1028 3145 1031
rect 3210 1028 3230 1031
rect 3234 1028 3262 1031
rect 3370 1028 3470 1031
rect 130 1018 134 1021
rect 194 1018 694 1021
rect 702 1018 710 1021
rect 714 1018 742 1021
rect 758 1021 761 1028
rect 758 1018 798 1021
rect 886 1018 894 1021
rect 910 1021 913 1028
rect 974 1022 977 1028
rect 3142 1022 3145 1028
rect 898 1018 913 1021
rect 938 1018 966 1021
rect 1018 1018 1094 1021
rect 1106 1018 1174 1021
rect 1186 1018 1198 1021
rect 1314 1018 1382 1021
rect 1450 1018 1462 1021
rect 1498 1018 1558 1021
rect 1674 1018 1950 1021
rect 1954 1018 1990 1021
rect 2026 1018 2478 1021
rect 2482 1018 2974 1021
rect 3058 1018 3078 1021
rect 90 1008 134 1011
rect 138 1008 326 1011
rect 530 1008 678 1011
rect 742 1011 745 1018
rect 1390 1012 1393 1018
rect 742 1008 822 1011
rect 866 1008 894 1011
rect 906 1008 1038 1011
rect 1066 1008 1102 1011
rect 1106 1008 1318 1011
rect 1402 1008 1486 1011
rect 1498 1008 1502 1011
rect 1602 1008 1670 1011
rect 1722 1008 1734 1011
rect 1746 1008 1790 1011
rect 1874 1008 1894 1011
rect 1898 1008 1934 1011
rect 1938 1008 2118 1011
rect 2122 1008 2270 1011
rect 2282 1008 2286 1011
rect 2298 1008 2342 1011
rect 2346 1008 2406 1011
rect 2706 1008 2718 1011
rect 2722 1008 2822 1011
rect 2850 1008 2942 1011
rect 2954 1008 2958 1011
rect 2978 1008 3182 1011
rect 3274 1008 3414 1011
rect 480 1003 482 1007
rect 486 1003 489 1007
rect 494 1003 496 1007
rect 1334 1002 1337 1008
rect 1512 1003 1514 1007
rect 1518 1003 1521 1007
rect 1526 1003 1528 1007
rect 1686 1002 1689 1008
rect 2536 1003 2538 1007
rect 2542 1003 2545 1007
rect 2550 1003 2552 1007
rect 714 998 734 1001
rect 786 998 902 1001
rect 946 998 958 1001
rect 970 998 974 1001
rect 1018 998 1046 1001
rect 1066 998 1086 1001
rect 1186 998 1326 1001
rect 1442 998 1470 1001
rect 1562 998 1598 1001
rect 1618 998 1678 1001
rect 1738 998 1902 1001
rect 1914 998 2006 1001
rect 2066 998 2070 1001
rect 2146 998 2206 1001
rect 2274 998 2486 1001
rect 2834 998 3014 1001
rect 3202 998 3510 1001
rect 3590 1001 3594 1002
rect 3562 998 3594 1001
rect 3526 992 3529 998
rect 302 988 366 991
rect 370 988 382 991
rect 458 988 534 991
rect 690 988 734 991
rect 874 988 910 991
rect 958 988 966 991
rect 970 988 998 991
rect 1010 988 1054 991
rect 1058 988 1086 991
rect 1138 988 1190 991
rect 1210 988 1214 991
rect 1250 988 1262 991
rect 1274 988 1358 991
rect 1370 988 1406 991
rect 1450 988 1534 991
rect 1586 988 1742 991
rect 1914 988 1982 991
rect 1986 988 2238 991
rect 2246 988 2254 991
rect 2258 988 2390 991
rect 2426 988 2430 991
rect 2642 988 3046 991
rect 3050 988 3134 991
rect 3138 988 3166 991
rect 302 982 305 988
rect 362 978 470 981
rect 514 978 694 981
rect 698 978 742 981
rect 818 978 1014 981
rect 1042 978 1078 981
rect 1082 978 1126 981
rect 1178 978 1305 981
rect 1314 978 1454 981
rect 1482 978 1918 981
rect 1922 978 2102 981
rect 2106 978 2286 981
rect 2290 978 2598 981
rect 2610 978 2614 981
rect 2618 978 2750 981
rect 2922 978 2926 981
rect 2930 978 2942 981
rect 2970 978 3110 981
rect 3422 981 3425 988
rect 3242 978 3425 981
rect 3590 981 3594 982
rect 3514 978 3594 981
rect 10 968 38 971
rect 242 968 286 971
rect 290 968 310 971
rect 442 968 1054 971
rect 1066 968 1118 971
rect 1154 968 1166 971
rect 1186 968 1230 971
rect 1302 971 1305 978
rect 1266 968 1289 971
rect 1302 968 1398 971
rect 1410 968 1414 971
rect 1418 968 1553 971
rect 1562 968 1582 971
rect 1586 968 1590 971
rect 1610 968 1646 971
rect 1674 968 1870 971
rect 1890 968 1950 971
rect 1962 968 2046 971
rect 2090 968 2110 971
rect 2174 968 2182 971
rect 2186 968 2190 971
rect 2194 968 2222 971
rect 2234 968 2238 971
rect 2242 968 2262 971
rect 2338 968 2350 971
rect 2362 968 2553 971
rect 2562 968 2894 971
rect 2906 968 3302 971
rect 3346 968 3350 971
rect 3378 968 3390 971
rect 3410 968 3542 971
rect 86 962 89 968
rect -26 961 -22 962
rect -26 958 6 961
rect 102 961 105 968
rect 158 961 161 968
rect 102 958 161 961
rect 298 958 382 961
rect 386 958 574 961
rect 578 958 630 961
rect 794 958 798 961
rect 834 958 1102 961
rect 1114 958 1126 961
rect 1146 958 1262 961
rect 1286 961 1289 968
rect 1286 958 1398 961
rect 1550 961 1553 968
rect 1550 958 1646 961
rect 1650 958 1718 961
rect 1754 958 1758 961
rect 1786 958 1798 961
rect 1810 958 1982 961
rect 2002 958 2014 961
rect 2174 961 2177 968
rect 2018 958 2177 961
rect 2186 958 2190 961
rect 2210 958 2366 961
rect 2370 958 2382 961
rect 2550 961 2553 968
rect 2550 958 2766 961
rect 2778 958 2801 961
rect 2810 958 2854 961
rect 2926 958 2958 961
rect 3154 958 3190 961
rect 3346 958 3433 961
rect 3466 958 3470 961
rect 694 952 697 958
rect 82 948 110 951
rect 186 948 222 951
rect 250 948 278 951
rect 290 948 329 951
rect 338 948 390 951
rect 394 948 414 951
rect 538 948 550 951
rect 610 948 646 951
rect 682 948 694 951
rect 762 948 782 951
rect 786 948 806 951
rect 858 948 878 951
rect 914 948 918 951
rect 954 948 982 951
rect 986 948 1006 951
rect 1050 948 1081 951
rect 1090 948 1134 951
rect 1154 948 1158 951
rect 1210 948 1214 951
rect 1226 948 1230 951
rect 1270 951 1273 958
rect 1270 948 1334 951
rect 1402 948 1470 951
rect 1514 948 1518 951
rect 1542 951 1545 958
rect 1542 948 1574 951
rect 1578 948 1582 951
rect 1610 948 1662 951
rect 1698 948 1742 951
rect 1746 948 1806 951
rect 1874 948 1878 951
rect 1898 948 1902 951
rect 1914 948 1966 951
rect 1970 948 1974 951
rect 1978 948 1990 951
rect 2026 948 2030 951
rect 2034 948 2158 951
rect 2186 948 2198 951
rect 2226 948 2326 951
rect 2330 948 2366 951
rect 2394 948 2446 951
rect 2546 948 2598 951
rect 2602 948 2654 951
rect 2730 948 2782 951
rect 2798 951 2801 958
rect 2926 952 2929 958
rect 2798 948 2926 951
rect 2938 948 2974 951
rect 2978 948 2982 951
rect 3086 951 3089 958
rect 3430 952 3433 958
rect 3074 948 3089 951
rect 3098 948 3102 951
rect 3146 948 3177 951
rect 3210 948 3214 951
rect 3242 948 3382 951
rect 3394 948 3422 951
rect 3434 948 3526 951
rect 34 938 70 941
rect 186 938 190 941
rect 258 938 318 941
rect 326 941 329 948
rect 326 938 358 941
rect 370 938 422 941
rect 474 938 526 941
rect 554 938 614 941
rect 730 938 750 941
rect 778 938 782 941
rect 790 938 846 941
rect 858 938 862 941
rect 986 938 990 941
rect 1042 938 1046 941
rect 1078 941 1081 948
rect 1254 942 1257 948
rect 1262 942 1265 948
rect 1678 942 1681 948
rect 2374 942 2377 948
rect 1078 938 1198 941
rect 1282 938 1318 941
rect 1418 938 1422 941
rect 1458 938 1465 941
rect 1474 938 1598 941
rect 1610 938 1630 941
rect 1722 938 1782 941
rect 1794 938 1798 941
rect 1810 938 1814 941
rect 1818 938 1846 941
rect 1858 938 1926 941
rect 1930 938 2054 941
rect 2066 938 2070 941
rect 2074 938 2118 941
rect 2154 938 2166 941
rect 2186 938 2198 941
rect 2226 938 2262 941
rect 2330 938 2334 941
rect 2418 938 2438 941
rect 2442 938 2462 941
rect 2662 941 2665 948
rect 2662 938 2774 941
rect 2834 938 2894 941
rect 2974 938 2982 941
rect 2998 941 3001 948
rect 3174 942 3177 948
rect 2986 938 3001 941
rect 3058 938 3078 941
rect 3194 938 3214 941
rect 3230 938 3233 948
rect 3242 938 3246 941
rect 3274 938 3278 941
rect 3314 938 3446 941
rect 170 928 182 931
rect 210 928 254 931
rect 282 928 398 931
rect 542 931 545 938
rect 790 932 793 938
rect 870 932 873 938
rect 910 932 913 938
rect 1054 932 1057 938
rect 1350 932 1353 938
rect 1462 932 1465 938
rect 1686 932 1689 938
rect 490 928 566 931
rect 606 928 614 931
rect 618 928 646 931
rect 650 928 782 931
rect 946 928 1030 931
rect 1098 928 1177 931
rect 1186 928 1238 931
rect 1282 928 1286 931
rect 1298 928 1302 931
rect 1306 928 1334 931
rect 1378 928 1390 931
rect 1394 928 1398 931
rect 1418 928 1446 931
rect 1482 928 1561 931
rect 1594 928 1670 931
rect 1730 928 1822 931
rect 1842 928 2046 931
rect 2090 928 2094 931
rect 2138 928 2390 931
rect 2714 928 2742 931
rect 2850 928 2918 931
rect 2970 928 3054 931
rect 3074 928 3078 931
rect 3130 928 3166 931
rect 3170 928 3222 931
rect 3250 928 3350 931
rect 3378 928 3406 931
rect 178 918 230 921
rect 270 921 273 928
rect 606 922 609 928
rect 270 918 294 921
rect 314 918 601 921
rect 634 918 726 921
rect 778 918 830 921
rect 882 918 926 921
rect 986 918 1038 921
rect 1050 918 1166 921
rect 1174 921 1177 928
rect 1174 918 1206 921
rect 1226 918 1342 921
rect 1362 918 1454 921
rect 1486 918 1494 921
rect 1498 918 1550 921
rect 1558 921 1561 928
rect 2062 922 2065 928
rect 1558 918 1710 921
rect 1722 918 1750 921
rect 1946 918 1950 921
rect 1978 918 2054 921
rect 2098 918 2102 921
rect 2298 918 2310 921
rect 2314 918 2510 921
rect 2742 921 2745 928
rect 2742 918 2798 921
rect 2950 921 2953 928
rect 2950 918 3102 921
rect 3122 918 3166 921
rect 3386 918 3406 921
rect 50 908 142 911
rect 258 908 422 911
rect 426 908 542 911
rect 598 911 601 918
rect 1918 912 1921 918
rect 1934 912 1937 918
rect 2710 912 2713 918
rect 598 908 670 911
rect 674 908 950 911
rect 970 908 982 911
rect 1026 908 1078 911
rect 1098 908 1230 911
rect 1242 908 1254 911
rect 1298 908 1302 911
rect 1322 908 1358 911
rect 1370 908 1406 911
rect 1418 908 1438 911
rect 1466 908 1518 911
rect 1522 908 1574 911
rect 1706 908 1798 911
rect 1810 908 1838 911
rect 1890 908 1894 911
rect 2050 908 2177 911
rect 2234 908 2302 911
rect 2306 908 2361 911
rect 2370 908 2638 911
rect 2722 908 2742 911
rect 2778 908 2862 911
rect 2882 908 2894 911
rect 2898 908 2982 911
rect 3106 908 3254 911
rect 3590 911 3594 912
rect 3394 908 3594 911
rect 992 903 994 907
rect 998 903 1001 907
rect 1006 903 1008 907
rect 2024 903 2026 907
rect 2030 903 2033 907
rect 2038 903 2040 907
rect 2174 902 2177 908
rect 218 898 294 901
rect 434 898 478 901
rect 562 898 782 901
rect 794 898 798 901
rect 866 898 926 901
rect 946 898 982 901
rect 1034 898 1214 901
rect 1250 898 1286 901
rect 1290 898 1302 901
rect 1306 898 1398 901
rect 1402 898 1486 901
rect 1490 898 1590 901
rect 1618 898 2017 901
rect 2138 898 2150 901
rect 2178 898 2198 901
rect 2346 898 2350 901
rect 2358 901 2361 908
rect 3040 903 3042 907
rect 3046 903 3049 907
rect 3054 903 3056 907
rect 2358 898 2382 901
rect 2698 898 2958 901
rect 2962 898 2974 901
rect 342 888 350 891
rect 354 888 462 891
rect 482 888 598 891
rect 634 888 790 891
rect 810 888 822 891
rect 842 888 854 891
rect 882 888 918 891
rect 938 888 990 891
rect 1002 888 1038 891
rect 1042 888 1054 891
rect 1114 888 1118 891
rect 1162 888 1174 891
rect 1210 888 1238 891
rect 1258 888 1270 891
rect 1282 888 1470 891
rect 1482 888 1550 891
rect 1562 888 1606 891
rect 1626 888 1654 891
rect 1670 888 1742 891
rect 1754 888 1846 891
rect 1850 888 1942 891
rect 1954 888 1958 891
rect 1986 888 2006 891
rect 2014 891 2017 898
rect 2014 888 2046 891
rect 2106 888 2134 891
rect 2190 888 2198 891
rect 2202 888 2262 891
rect 2282 888 2390 891
rect 2434 888 2457 891
rect 2466 888 2614 891
rect 2626 888 2758 891
rect 2790 888 2814 891
rect 2826 888 2942 891
rect 2946 888 2966 891
rect 2994 888 3030 891
rect 3034 888 3038 891
rect 3042 888 3046 891
rect 3102 888 3206 891
rect 3590 891 3594 892
rect 3346 888 3594 891
rect 18 878 30 881
rect 58 878 62 881
rect 286 881 289 888
rect 286 878 326 881
rect 330 878 366 881
rect 370 878 398 881
rect 410 878 454 881
rect 490 878 518 881
rect 538 878 622 881
rect 634 878 702 881
rect 722 878 798 881
rect 802 878 806 881
rect 834 878 910 881
rect 962 878 998 881
rect 1026 878 1062 881
rect 1074 878 1150 881
rect 1162 878 1166 881
rect 1246 881 1249 888
rect 1670 882 1673 888
rect 2454 882 2457 888
rect 2790 882 2793 888
rect 3102 882 3105 888
rect 1194 878 1233 881
rect 1246 878 1270 881
rect 1282 878 1350 881
rect 1370 878 1478 881
rect 1498 878 1614 881
rect 1626 878 1646 881
rect 1682 878 1694 881
rect 1706 878 1766 881
rect 1802 878 1958 881
rect 1978 878 2230 881
rect 2466 878 2470 881
rect 2746 878 2750 881
rect 2770 878 2790 881
rect 2802 878 2854 881
rect 2906 878 2926 881
rect 2986 878 3030 881
rect 3034 878 3054 881
rect 3058 878 3078 881
rect 3170 878 3222 881
rect 3226 878 3278 881
rect 3282 878 3334 881
rect 3338 878 3390 881
rect 18 868 78 871
rect 114 868 206 871
rect 254 871 257 878
rect 1230 872 1233 878
rect 1702 872 1705 878
rect 2302 872 2305 878
rect 2310 872 2313 878
rect 226 868 257 871
rect 322 868 430 871
rect 474 868 502 871
rect 562 868 582 871
rect 618 868 686 871
rect 698 868 742 871
rect 778 868 902 871
rect 994 868 1030 871
rect 1106 868 1174 871
rect 1186 868 1198 871
rect 1242 868 1310 871
rect 1330 868 1334 871
rect 1346 868 1422 871
rect 1434 868 1486 871
rect 1538 868 1582 871
rect 1610 868 1697 871
rect 1754 868 1814 871
rect 1826 868 2038 871
rect 2058 868 2070 871
rect 2090 868 2113 871
rect 2122 868 2126 871
rect 2154 868 2158 871
rect 2202 868 2206 871
rect 2250 868 2270 871
rect 2350 871 2353 878
rect 2314 868 2353 871
rect 2446 872 2449 878
rect 2518 872 2521 878
rect 2506 868 2510 871
rect 2610 868 2614 871
rect 2682 868 3494 871
rect 3518 868 3526 871
rect 3590 871 3594 872
rect 3530 868 3594 871
rect 614 862 617 868
rect 950 862 953 868
rect 82 858 94 861
rect 98 858 134 861
rect 138 858 166 861
rect 202 858 214 861
rect 234 858 238 861
rect 242 858 286 861
rect 314 858 334 861
rect 346 858 350 861
rect 450 858 550 861
rect 634 858 718 861
rect 730 858 758 861
rect 802 858 806 861
rect 834 858 838 861
rect 858 858 862 861
rect 874 858 878 861
rect 978 858 1014 861
rect 1018 858 1062 861
rect 1082 858 1094 861
rect 1146 858 1310 861
rect 1322 858 1326 861
rect 1338 858 1342 861
rect 1386 858 1390 861
rect 1402 858 1558 861
rect 1570 858 1574 861
rect 1578 858 1590 861
rect 1666 858 1670 861
rect 1694 861 1697 868
rect 1694 858 1726 861
rect 1738 858 1758 861
rect 1762 858 1774 861
rect 1834 858 1894 861
rect 1938 858 1942 861
rect 1962 858 1982 861
rect 1986 858 1990 861
rect 1994 858 2070 861
rect 2074 858 2102 861
rect 2110 861 2113 868
rect 2110 858 2142 861
rect 2154 858 2342 861
rect 2410 858 2414 861
rect 2434 858 2438 861
rect 2442 858 2494 861
rect 2586 858 2678 861
rect 2682 858 2686 861
rect 2786 858 2838 861
rect 2866 858 2870 861
rect 2906 858 2926 861
rect 2938 858 3286 861
rect 3290 858 3342 861
rect 3410 858 3414 861
rect 622 852 625 858
rect 1118 852 1121 858
rect 66 848 110 851
rect 130 848 182 851
rect 290 848 510 851
rect 674 848 686 851
rect 702 848 814 851
rect 818 848 878 851
rect 986 848 1110 851
rect 1130 848 1150 851
rect 1178 848 1198 851
rect 1210 848 1294 851
rect 1386 848 1390 851
rect 1410 848 1414 851
rect 1426 848 1430 851
rect 1450 848 1462 851
rect 1474 848 1478 851
rect 1554 848 1574 851
rect 1582 848 1590 851
rect 1594 848 1662 851
rect 1678 851 1681 858
rect 1674 848 1681 851
rect 1690 848 1822 851
rect 1842 848 1886 851
rect 1930 848 1934 851
rect 1962 848 1966 851
rect 2050 848 2054 851
rect 2082 848 2086 851
rect 2110 848 2126 851
rect 2234 848 2238 851
rect 2378 848 2486 851
rect 2506 848 2518 851
rect 2658 848 2678 851
rect 2694 848 2878 851
rect 2914 848 2985 851
rect 2994 848 3086 851
rect 3106 848 3126 851
rect 3138 848 3174 851
rect 3226 848 3230 851
rect 3426 848 3526 851
rect 3590 851 3594 852
rect 3562 848 3594 851
rect 54 841 57 848
rect 518 842 521 848
rect 582 842 585 848
rect 702 842 705 848
rect 966 842 969 848
rect 54 838 70 841
rect 90 838 118 841
rect 130 838 190 841
rect 266 838 446 841
rect 458 838 494 841
rect 682 838 702 841
rect 722 838 726 841
rect 754 838 846 841
rect 922 838 950 841
rect 978 838 1046 841
rect 1058 838 1254 841
rect 1306 838 1358 841
rect 1378 838 1438 841
rect 1450 838 1454 841
rect 1482 838 1494 841
rect 1554 838 1766 841
rect 1770 838 1910 841
rect 1934 841 1937 848
rect 2110 842 2113 848
rect 2294 842 2297 848
rect 1934 838 1982 841
rect 2042 838 2070 841
rect 2138 838 2158 841
rect 2162 838 2262 841
rect 2326 841 2329 848
rect 2694 842 2697 848
rect 2326 838 2470 841
rect 2674 838 2694 841
rect 2714 838 2774 841
rect 2778 838 2934 841
rect 2982 841 2985 848
rect 2982 838 2998 841
rect 3018 838 3118 841
rect 3130 838 3166 841
rect 58 828 62 831
rect 178 828 526 831
rect 590 831 593 838
rect 598 831 601 838
rect 590 828 601 831
rect 614 831 617 838
rect 610 828 617 831
rect 642 828 662 831
rect 666 828 766 831
rect 778 828 822 831
rect 850 828 926 831
rect 930 828 1038 831
rect 1050 828 1054 831
rect 1114 828 1126 831
rect 1202 828 1222 831
rect 1242 828 1246 831
rect 1258 828 1550 831
rect 1562 828 1566 831
rect 1578 828 1606 831
rect 1618 828 1630 831
rect 1638 828 1646 831
rect 1650 828 1806 831
rect 2590 831 2593 838
rect 1814 828 3062 831
rect 3590 831 3594 832
rect 3498 828 3594 831
rect 242 818 334 821
rect 354 818 406 821
rect 410 818 505 821
rect 570 818 598 821
rect 1814 821 1817 828
rect 618 818 1817 821
rect 1898 818 1902 821
rect 1926 818 2022 821
rect 2042 818 2286 821
rect 2450 818 2550 821
rect 2650 818 2678 821
rect 2706 818 2710 821
rect 2714 818 2750 821
rect 2754 818 2806 821
rect 2810 818 2830 821
rect 2890 818 3254 821
rect 50 808 126 811
rect 130 808 206 811
rect 210 808 334 811
rect 354 808 358 811
rect 426 808 462 811
rect 502 811 505 818
rect 502 808 790 811
rect 810 808 886 811
rect 906 808 974 811
rect 986 808 990 811
rect 1002 808 1182 811
rect 1210 808 1262 811
rect 1298 808 1342 811
rect 1370 808 1382 811
rect 1394 808 1398 811
rect 1410 808 1462 811
rect 1546 808 1654 811
rect 1706 808 1718 811
rect 1926 811 1929 818
rect 1762 808 1929 811
rect 1938 808 2094 811
rect 2114 808 2254 811
rect 2682 808 2950 811
rect 3082 808 3094 811
rect 3590 811 3594 812
rect 3474 808 3594 811
rect 480 803 482 807
rect 486 803 489 807
rect 494 803 496 807
rect 1512 803 1514 807
rect 1518 803 1521 807
rect 1526 803 1528 807
rect 2536 803 2538 807
rect 2542 803 2545 807
rect 2550 803 2552 807
rect 154 798 182 801
rect 186 798 270 801
rect 402 798 454 801
rect 458 798 470 801
rect 594 798 630 801
rect 730 798 766 801
rect 786 798 790 801
rect 818 798 886 801
rect 890 798 982 801
rect 1074 798 1246 801
rect 1258 798 1302 801
rect 1314 798 1318 801
rect 1362 798 1494 801
rect 1658 798 1750 801
rect 1802 798 1878 801
rect 1882 798 1902 801
rect 1914 798 1950 801
rect 2154 798 2390 801
rect 2410 798 2526 801
rect 2570 798 2782 801
rect 2786 798 3134 801
rect 3378 798 3398 801
rect 1638 792 1641 798
rect 186 788 678 791
rect 742 788 958 791
rect 994 788 1166 791
rect 1202 788 1222 791
rect 1226 788 1334 791
rect 1354 788 1374 791
rect 1394 788 1478 791
rect 1506 788 1510 791
rect 1530 788 1542 791
rect 1674 788 1694 791
rect 1714 788 1798 791
rect 1834 788 1902 791
rect 1914 788 1942 791
rect 2002 788 2014 791
rect 2210 788 2406 791
rect 2426 788 2438 791
rect 2490 788 2598 791
rect 2610 788 2798 791
rect 2802 788 3502 791
rect 3590 791 3594 792
rect 3562 788 3594 791
rect 338 778 502 781
rect 734 781 737 788
rect 582 778 737 781
rect 742 782 745 788
rect 786 778 822 781
rect 834 778 1150 781
rect 1162 778 1238 781
rect 1314 778 1334 781
rect 1434 778 2566 781
rect 2634 778 2646 781
rect 2858 778 2902 781
rect 2962 778 2966 781
rect 2970 778 3214 781
rect 3466 778 3478 781
rect 3518 781 3521 788
rect 3518 778 3593 781
rect 582 772 585 778
rect 210 768 246 771
rect 466 768 566 771
rect 722 768 758 771
rect 762 768 814 771
rect 882 768 918 771
rect 938 768 1118 771
rect 1122 768 1134 771
rect 1146 768 1174 771
rect 1178 768 1206 771
rect 1246 771 1249 778
rect 1342 771 1345 778
rect 3590 772 3593 778
rect 1246 768 1345 771
rect 1354 768 1390 771
rect 1418 768 1486 771
rect 1566 768 1574 771
rect 1610 768 1614 771
rect 1634 768 1638 771
rect 1658 768 1774 771
rect 1818 768 2046 771
rect 2058 768 2062 771
rect 2070 768 2094 771
rect 2114 768 2630 771
rect 2738 768 2742 771
rect 2786 768 3086 771
rect 3106 768 3142 771
rect 3182 768 3262 771
rect 3538 768 3550 771
rect 3590 768 3594 772
rect 262 761 265 768
rect 234 758 265 761
rect 298 758 302 761
rect 318 761 321 768
rect 318 758 366 761
rect 370 758 390 761
rect 426 758 438 761
rect 566 761 569 768
rect 566 758 710 761
rect 722 758 822 761
rect 826 758 838 761
rect 858 758 894 761
rect 926 761 929 768
rect 1230 762 1233 768
rect 906 758 929 761
rect 1002 758 1006 761
rect 1066 758 1070 761
rect 1146 758 1206 761
rect 1242 758 1270 761
rect 1290 758 1350 761
rect 1450 758 1590 761
rect 1814 761 1817 768
rect 2070 762 2073 768
rect 3182 762 3185 768
rect 1602 758 1817 761
rect 1834 758 1942 761
rect 1986 758 1990 761
rect 1994 758 2046 761
rect 2078 758 2150 761
rect 2154 758 2158 761
rect 2170 758 2222 761
rect 2298 758 2334 761
rect 2410 758 2414 761
rect 2422 758 2430 761
rect 2434 758 2446 761
rect 2642 758 3094 761
rect 3162 758 3166 761
rect 3218 758 3478 761
rect 82 748 278 751
rect 362 748 390 751
rect 394 748 462 751
rect 466 748 478 751
rect 482 748 518 751
rect 522 748 550 751
rect 554 748 574 751
rect 610 748 625 751
rect 650 748 721 751
rect 730 748 846 751
rect 858 748 1590 751
rect 1626 748 1662 751
rect 1686 748 1726 751
rect 1834 748 1838 751
rect 1882 748 1998 751
rect 2078 751 2081 758
rect 2034 748 2081 751
rect 2090 748 2118 751
rect 2130 748 2134 751
rect 2162 748 2174 751
rect 2194 748 2198 751
rect 2282 748 2286 751
rect 2342 751 2345 758
rect 2314 748 2345 751
rect 2410 748 2438 751
rect 2534 751 2537 758
rect 2506 748 2537 751
rect 2570 748 2622 751
rect 2714 748 2758 751
rect 2762 748 2766 751
rect 2778 748 2838 751
rect 2850 748 2894 751
rect 582 742 585 748
rect 622 742 625 748
rect 50 738 62 741
rect 98 738 110 741
rect 258 738 302 741
rect 322 738 374 741
rect 378 738 510 741
rect 514 738 542 741
rect 570 738 574 741
rect 674 738 702 741
rect 718 741 721 748
rect 1686 742 1689 748
rect 1734 742 1737 748
rect 1862 742 1865 748
rect 2470 742 2473 748
rect 718 738 742 741
rect 746 738 766 741
rect 882 738 886 741
rect 890 738 982 741
rect 1054 738 1062 741
rect 1066 738 1078 741
rect 1082 738 1126 741
rect 1146 738 1166 741
rect 1186 738 1198 741
rect 1210 738 1286 741
rect 1306 738 1310 741
rect 1330 738 1334 741
rect 1346 738 1350 741
rect 1418 738 1422 741
rect 1434 738 1545 741
rect 1554 738 1582 741
rect 1594 738 1654 741
rect 1714 738 1726 741
rect 1754 738 1782 741
rect 1786 738 1830 741
rect 1834 738 1838 741
rect 1866 738 1894 741
rect 1954 738 1958 741
rect 1994 738 2006 741
rect 2026 738 2214 741
rect 2226 738 2230 741
rect 2250 738 2270 741
rect 2290 738 2462 741
rect 2550 741 2553 748
rect 2906 748 2961 751
rect 2958 742 2961 748
rect 3042 748 3062 751
rect 3102 751 3105 758
rect 3102 748 3190 751
rect 3194 748 3222 751
rect 3290 748 3438 751
rect 3590 751 3594 752
rect 3450 748 3594 751
rect 2974 742 2977 748
rect 3390 742 3393 748
rect 2550 738 2614 741
rect 2626 738 2654 741
rect 2658 738 2726 741
rect 2746 738 2750 741
rect 2770 738 2790 741
rect 3002 738 3006 741
rect 3034 738 3078 741
rect 3098 738 3118 741
rect 3202 738 3294 741
rect 182 732 185 738
rect 558 732 561 738
rect 814 732 817 738
rect 1030 732 1033 738
rect 50 728 54 731
rect 74 728 86 731
rect 90 728 174 731
rect 306 728 374 731
rect 434 728 462 731
rect 586 728 662 731
rect 666 728 694 731
rect 714 728 734 731
rect 874 728 886 731
rect 946 728 950 731
rect 970 728 974 731
rect 1142 731 1145 738
rect 1098 728 1145 731
rect 1154 728 1230 731
rect 1242 728 1246 731
rect 1258 728 1310 731
rect 1330 728 1374 731
rect 1406 728 1409 738
rect 1542 732 1545 738
rect 2726 732 2729 738
rect 1482 728 1510 731
rect 1546 728 1582 731
rect 1586 728 1670 731
rect 1722 728 1742 731
rect 1746 728 1766 731
rect 1786 728 1934 731
rect 1954 728 1958 731
rect 2006 728 2014 731
rect 2018 728 2054 731
rect 2094 728 2102 731
rect 2106 728 2118 731
rect 2130 728 2318 731
rect 2418 728 2422 731
rect 2458 728 2478 731
rect 2498 728 2606 731
rect 2626 728 2630 731
rect 2658 728 2662 731
rect 2730 728 2822 731
rect 2826 728 2854 731
rect 2962 728 3038 731
rect 3042 728 3054 731
rect 3178 728 3222 731
rect 3234 728 3326 731
rect 3330 728 3430 731
rect 414 722 417 728
rect 122 718 142 721
rect 274 718 350 721
rect 466 718 542 721
rect 562 718 638 721
rect 658 718 870 721
rect 882 718 998 721
rect 1042 718 1070 721
rect 1074 718 1102 721
rect 1106 718 1126 721
rect 1138 718 1454 721
rect 1470 721 1473 728
rect 1470 718 1486 721
rect 1498 718 1502 721
rect 1594 718 1614 721
rect 1626 718 1654 721
rect 1726 718 1734 721
rect 1738 718 1854 721
rect 1866 718 1934 721
rect 1974 721 1977 728
rect 1974 718 1998 721
rect 2002 718 2054 721
rect 2062 721 2065 728
rect 2062 718 2134 721
rect 2162 718 2174 721
rect 2282 718 2286 721
rect 2370 718 2398 721
rect 2618 718 2742 721
rect 2794 718 2806 721
rect 2866 718 2870 721
rect 2878 718 3198 721
rect 3202 718 3454 721
rect 1566 712 1569 718
rect 34 708 38 711
rect 186 708 262 711
rect 266 708 438 711
rect 474 708 878 711
rect 962 708 974 711
rect 1034 708 1110 711
rect 1162 708 1166 711
rect 1178 708 1182 711
rect 1290 708 1294 711
rect 1442 708 1446 711
rect 1482 708 1558 711
rect 1650 708 1830 711
rect 1946 708 2014 711
rect 2106 708 2262 711
rect 2314 708 2334 711
rect 2346 708 2374 711
rect 2378 708 2542 711
rect 2562 708 2566 711
rect 2738 708 2806 711
rect 2878 711 2881 718
rect 2810 708 2881 711
rect 2890 708 2894 711
rect 2962 708 2982 711
rect 3002 708 3030 711
rect 3114 708 3142 711
rect 3162 708 3198 711
rect 3338 708 3422 711
rect 886 702 889 708
rect 992 703 994 707
rect 998 703 1001 707
rect 1006 703 1008 707
rect 2024 703 2026 707
rect 2030 703 2033 707
rect 2038 703 2040 707
rect 3040 703 3042 707
rect 3046 703 3049 707
rect 3054 703 3056 707
rect 26 698 158 701
rect 162 698 206 701
rect 210 698 246 701
rect 258 698 590 701
rect 626 698 718 701
rect 730 698 742 701
rect 746 698 766 701
rect 786 698 878 701
rect 962 698 982 701
rect 1042 698 1190 701
rect 1194 698 1230 701
rect 1242 698 1398 701
rect 1402 698 1622 701
rect 1650 698 1790 701
rect 1802 698 1822 701
rect 1826 698 2014 701
rect 2178 698 2366 701
rect 2394 698 2814 701
rect 2858 698 2910 701
rect 2914 698 2990 701
rect 3226 698 3358 701
rect 726 692 729 698
rect 3206 692 3209 698
rect 190 688 310 691
rect 506 688 606 691
rect 610 688 718 691
rect 754 688 774 691
rect 914 688 918 691
rect 930 688 1038 691
rect 1138 688 1158 691
rect 1210 688 1318 691
rect 1470 688 1582 691
rect 1590 688 1678 691
rect 1682 688 1710 691
rect 1718 688 1726 691
rect 1730 688 1734 691
rect 1762 688 1774 691
rect 1818 688 1822 691
rect 1834 688 1846 691
rect 1858 688 1870 691
rect 1890 688 2166 691
rect 2226 688 2318 691
rect 2322 688 2326 691
rect 2330 688 2350 691
rect 2402 688 2494 691
rect 2602 688 2654 691
rect 2762 688 2926 691
rect 2930 688 2990 691
rect 3018 688 3110 691
rect 3154 688 3158 691
rect 3218 688 3310 691
rect 3426 688 3510 691
rect 3514 688 3526 691
rect 190 682 193 688
rect 18 678 38 681
rect 74 678 110 681
rect 114 678 182 681
rect 322 678 366 681
rect 370 678 414 681
rect 418 678 470 681
rect 490 678 518 681
rect 522 678 526 681
rect 546 678 726 681
rect 862 678 870 681
rect 874 678 966 681
rect 986 678 1070 681
rect 1078 681 1081 688
rect 1342 682 1345 688
rect 1470 682 1473 688
rect 1590 682 1593 688
rect 2398 682 2401 688
rect 1078 678 1086 681
rect 1122 678 1126 681
rect 1138 678 1142 681
rect 1154 678 1206 681
rect 1218 678 1230 681
rect 1242 678 1278 681
rect 1282 678 1310 681
rect 1330 678 1334 681
rect 1362 678 1366 681
rect 1370 678 1390 681
rect 1402 678 1430 681
rect 1506 678 1510 681
rect 1522 678 1590 681
rect 1610 678 1614 681
rect 1658 678 1662 681
rect 1722 678 1726 681
rect 1770 678 1910 681
rect 1914 678 1950 681
rect 2018 678 2070 681
rect 2130 678 2182 681
rect 2218 678 2310 681
rect 2314 678 2334 681
rect 2338 678 2398 681
rect 2410 678 2414 681
rect 2530 678 2622 681
rect 2662 681 2665 688
rect 2662 678 2694 681
rect 2710 681 2713 688
rect 2710 678 2726 681
rect 2746 678 2870 681
rect 3026 678 3038 681
rect 3082 678 3094 681
rect 3106 678 3110 681
rect 3114 678 3222 681
rect 3230 678 3366 681
rect 42 668 78 671
rect 122 668 126 671
rect 138 668 198 671
rect 282 668 334 671
rect 378 668 662 671
rect 666 668 670 671
rect 682 668 686 671
rect 738 668 806 671
rect 834 668 838 671
rect 982 671 985 678
rect 850 668 985 671
rect 1034 668 1262 671
rect 1290 668 1470 671
rect 1514 668 1694 671
rect 1706 668 1718 671
rect 1738 668 1769 671
rect 1778 668 1782 671
rect 1794 668 1886 671
rect 2006 671 2009 678
rect 1890 668 2009 671
rect 2018 668 2022 671
rect 2078 671 2081 678
rect 2438 672 2441 678
rect 2078 668 2110 671
rect 2194 668 2206 671
rect 2370 668 2374 671
rect 2410 668 2430 671
rect 2770 668 2878 671
rect 2954 668 2974 671
rect 3006 671 3009 678
rect 3006 668 3062 671
rect 3082 668 3118 671
rect 3154 668 3214 671
rect 3230 671 3233 678
rect 3226 668 3233 671
rect 3238 668 3326 671
rect 3366 671 3369 678
rect 3366 668 3414 671
rect 1766 662 1769 668
rect 2150 662 2153 668
rect 18 658 94 661
rect 98 658 142 661
rect 186 658 238 661
rect 338 658 342 661
rect 386 658 390 661
rect 450 658 454 661
rect 474 658 526 661
rect 562 658 590 661
rect 610 658 750 661
rect 794 658 870 661
rect 874 658 958 661
rect 962 658 1006 661
rect 1010 658 1222 661
rect 1234 658 1238 661
rect 1250 658 1254 661
rect 1274 658 1278 661
rect 1290 658 1294 661
rect 1322 658 1366 661
rect 1402 658 1406 661
rect 1466 658 1494 661
rect 1594 658 1614 661
rect 1618 658 1646 661
rect 1650 658 1758 661
rect 1850 658 1854 661
rect 1890 658 1910 661
rect 1930 658 2014 661
rect 2058 658 2062 661
rect 2082 658 2086 661
rect 2130 658 2134 661
rect 2286 661 2289 668
rect 2646 662 2649 668
rect 2218 658 2342 661
rect 2482 658 2561 661
rect 2678 661 2681 668
rect 2678 658 2742 661
rect 2746 658 2790 661
rect 2802 658 2814 661
rect 2890 658 2894 661
rect 2906 658 3070 661
rect 3074 658 3110 661
rect 3130 658 3166 661
rect 3186 658 3206 661
rect 3238 661 3241 668
rect 3210 658 3241 661
rect 3250 659 3262 661
rect 3250 658 3265 659
rect 3322 658 3518 661
rect 66 648 198 651
rect 258 648 262 651
rect 302 651 305 658
rect 298 648 305 651
rect 462 651 465 658
rect 394 648 465 651
rect 518 652 521 658
rect 594 648 646 651
rect 658 648 702 651
rect 714 648 718 651
rect 730 648 1366 651
rect 1378 648 1430 651
rect 1458 648 1462 651
rect 1482 648 1542 651
rect 1554 648 1662 651
rect 1690 648 1750 651
rect 1906 648 2046 651
rect 2070 648 2094 651
rect 2198 651 2201 658
rect 2558 652 2561 658
rect 2198 648 2254 651
rect 2330 648 2366 651
rect 2394 648 2462 651
rect 2690 648 2694 651
rect 2706 648 2742 651
rect 2838 651 2841 658
rect 2838 648 2921 651
rect 2930 648 3294 651
rect 3362 648 3454 651
rect 3590 651 3594 652
rect 3562 648 3594 651
rect 66 638 214 641
rect 218 638 270 641
rect 286 641 289 648
rect 382 642 385 648
rect 2070 642 2073 648
rect 286 638 382 641
rect 394 638 430 641
rect 514 638 534 641
rect 610 638 614 641
rect 682 638 694 641
rect 702 638 945 641
rect 954 638 958 641
rect 970 638 1054 641
rect 1058 638 1062 641
rect 90 628 150 631
rect 154 628 222 631
rect 234 628 398 631
rect 434 628 478 631
rect 702 631 705 638
rect 586 628 705 631
rect 714 628 894 631
rect 914 628 918 631
rect 942 631 945 638
rect 1070 632 1073 638
rect 942 628 1014 631
rect 1102 631 1105 638
rect 1198 631 1201 638
rect 1102 628 1201 631
rect 1206 632 1209 638
rect 1214 632 1217 641
rect 1274 638 1286 641
rect 1346 638 1422 641
rect 1434 638 1526 641
rect 1562 638 1734 641
rect 1822 638 1862 641
rect 1866 638 1870 641
rect 1890 638 1894 641
rect 1922 638 1926 641
rect 1938 638 1942 641
rect 2082 638 2086 641
rect 2130 638 2134 641
rect 2170 638 2286 641
rect 2386 638 2406 641
rect 2462 638 2470 641
rect 2474 638 2494 641
rect 2514 638 2630 641
rect 2634 638 2774 641
rect 2890 638 2902 641
rect 2918 641 2921 648
rect 2918 638 2990 641
rect 3042 638 3046 641
rect 3102 638 3134 641
rect 3194 638 3198 641
rect 3210 638 3214 641
rect 3370 638 3374 641
rect 3394 638 3526 641
rect 1226 628 1358 631
rect 1410 628 1462 631
rect 1490 628 1550 631
rect 1602 628 1614 631
rect 1682 628 1694 631
rect 1822 631 1825 638
rect 1698 628 1825 631
rect 2846 631 2849 638
rect 3102 632 3105 638
rect 1834 628 2849 631
rect 2926 628 2958 631
rect 414 622 417 628
rect 2926 622 2929 628
rect 154 618 374 621
rect 434 618 614 621
rect 698 618 1086 621
rect 1090 618 1094 621
rect 1178 618 1182 621
rect 1258 618 1358 621
rect 1506 618 1550 621
rect 1626 618 2174 621
rect 2482 618 2542 621
rect 2674 618 2710 621
rect 2938 618 2974 621
rect 3034 618 3342 621
rect 146 608 374 611
rect 562 608 662 611
rect 666 608 822 611
rect 874 608 1118 611
rect 1122 608 1238 611
rect 1274 608 1334 611
rect 1346 608 1374 611
rect 1578 608 1710 611
rect 1934 608 1942 611
rect 2378 608 2526 611
rect 2626 608 2998 611
rect 3026 608 3198 611
rect 480 603 482 607
rect 486 603 489 607
rect 494 603 496 607
rect 1512 603 1514 607
rect 1518 603 1521 607
rect 1526 603 1528 607
rect 1934 602 1937 608
rect 2536 603 2538 607
rect 2542 603 2545 607
rect 2550 603 2552 607
rect 186 598 470 601
rect 502 598 1414 601
rect 1554 598 1574 601
rect 1578 598 1822 601
rect 1826 598 1934 601
rect 1986 598 2110 601
rect 2562 598 2990 601
rect 3058 598 3110 601
rect 58 588 238 591
rect 502 591 505 598
rect 274 588 505 591
rect 578 588 654 591
rect 658 588 838 591
rect 878 588 886 591
rect 906 588 934 591
rect 946 588 1022 591
rect 1042 588 1046 591
rect 1058 588 2862 591
rect 3074 588 3286 591
rect 3290 588 3406 591
rect 154 578 278 581
rect 366 578 374 581
rect 378 578 582 581
rect 690 578 766 581
rect 778 578 790 581
rect 802 578 878 581
rect 882 578 1126 581
rect 1154 578 1190 581
rect 1202 578 1334 581
rect 1386 578 1558 581
rect 1610 578 1958 581
rect 1994 578 1998 581
rect 2114 578 2166 581
rect 2170 578 2206 581
rect 2322 578 2358 581
rect 2378 578 2422 581
rect 2434 578 2558 581
rect 2618 578 2654 581
rect 2866 578 2870 581
rect 3066 578 3102 581
rect 114 568 182 571
rect 334 571 337 578
rect 334 568 422 571
rect 642 568 694 571
rect 722 568 737 571
rect 754 568 766 571
rect 770 568 782 571
rect 810 568 910 571
rect 918 568 1198 571
rect 1314 568 1318 571
rect 1330 568 1502 571
rect 1506 568 1550 571
rect 1658 568 1734 571
rect 1754 568 1798 571
rect 1866 568 2286 571
rect 2290 568 2638 571
rect 2642 568 2870 571
rect 2962 568 3086 571
rect 3114 568 3142 571
rect 3534 568 3542 571
rect 3590 571 3594 572
rect 3546 568 3594 571
rect 734 562 737 568
rect 106 558 134 561
rect 138 558 166 561
rect 170 558 238 561
rect 242 558 286 561
rect 306 558 310 561
rect 498 558 502 561
rect 546 558 630 561
rect 698 558 710 561
rect 754 558 910 561
rect 918 561 921 568
rect 914 558 921 561
rect 938 558 958 561
rect 962 558 982 561
rect 1010 558 1073 561
rect 1086 558 1094 561
rect 1098 558 1102 561
rect 1118 558 1134 561
rect 1170 558 1222 561
rect 1226 558 1270 561
rect 1282 558 1286 561
rect 1294 561 1297 568
rect 1294 558 1366 561
rect 1426 558 1518 561
rect 1602 558 1694 561
rect 1746 558 1774 561
rect 1810 558 1814 561
rect 1842 558 1894 561
rect 1922 558 1998 561
rect 2046 558 2070 561
rect 2122 558 2150 561
rect 2162 558 2278 561
rect 2282 558 2342 561
rect 2358 558 2446 561
rect 2586 558 2598 561
rect 2650 558 2686 561
rect 2762 558 2774 561
rect 2782 558 2926 561
rect 2934 558 2966 561
rect 3002 558 3030 561
rect 3050 558 3094 561
rect 3106 558 3238 561
rect 6 548 14 551
rect 18 548 46 551
rect 70 551 73 558
rect 50 548 73 551
rect 114 548 190 551
rect 334 551 337 558
rect 926 552 929 558
rect 1070 552 1073 558
rect 1110 552 1113 558
rect 1118 552 1121 558
rect 1142 552 1145 558
rect 2046 552 2049 558
rect 194 548 337 551
rect 570 548 574 551
rect 610 548 662 551
rect 778 548 830 551
rect 850 548 854 551
rect 858 548 902 551
rect 946 548 1030 551
rect 1034 548 1062 551
rect 1130 548 1134 551
rect 1162 548 1198 551
rect 1250 548 1321 551
rect 1338 548 1345 551
rect 1386 548 1390 551
rect 1410 548 1417 551
rect 70 541 73 548
rect 70 538 214 541
rect 322 538 414 541
rect 518 541 521 548
rect 606 542 609 548
rect 518 538 598 541
rect 626 538 654 541
rect 742 541 745 548
rect 1318 542 1321 548
rect 1342 542 1345 548
rect 1414 542 1417 548
rect 1482 548 1486 551
rect 1594 548 1654 551
rect 1690 548 1729 551
rect 1738 548 1766 551
rect 1794 548 1870 551
rect 1906 548 1918 551
rect 1930 548 1977 551
rect 1994 548 1998 551
rect 2154 548 2201 551
rect 2358 551 2361 558
rect 2314 548 2361 551
rect 2370 548 2382 551
rect 2458 548 2510 551
rect 2582 548 2678 551
rect 2734 551 2737 558
rect 2722 548 2737 551
rect 2782 551 2785 558
rect 2746 548 2785 551
rect 2802 548 2806 551
rect 2934 551 2937 558
rect 2914 548 2937 551
rect 3002 548 3009 551
rect 3018 548 3070 551
rect 3162 548 3166 551
rect 3178 548 3182 551
rect 3202 548 3230 551
rect 3242 548 3278 551
rect 3422 551 3425 558
rect 3322 548 3425 551
rect 3590 551 3594 552
rect 3514 548 3594 551
rect 1454 542 1457 548
rect 738 538 745 541
rect 754 538 838 541
rect 842 538 886 541
rect 906 538 990 541
rect 1082 538 1086 541
rect 1138 538 1150 541
rect 1178 538 1182 541
rect 1194 538 1310 541
rect 1538 538 1598 541
rect 1642 538 1646 541
rect 1714 538 1718 541
rect 1726 541 1729 548
rect 1902 541 1905 548
rect 1726 538 1905 541
rect 1914 538 1950 541
rect 1962 538 1966 541
rect 1974 541 1977 548
rect 2198 542 2201 548
rect 2582 542 2585 548
rect 2678 542 2681 548
rect 1974 538 1998 541
rect 2010 538 2134 541
rect 2306 538 2358 541
rect 2506 538 2542 541
rect 2626 538 2670 541
rect 2690 538 2742 541
rect 2746 538 2806 541
rect 2890 538 2926 541
rect 2950 541 2953 548
rect 2982 541 2985 548
rect 3294 542 3297 548
rect 2946 538 2985 541
rect 3010 538 3014 541
rect 3042 538 3086 541
rect 3090 538 3230 541
rect 3298 538 3326 541
rect 3346 538 3486 541
rect 3490 538 3494 541
rect 1046 532 1049 538
rect 202 528 206 531
rect 226 528 358 531
rect 362 528 398 531
rect 410 528 414 531
rect 426 528 798 531
rect 874 528 926 531
rect 978 528 1014 531
rect 1066 528 1198 531
rect 1226 528 1438 531
rect 1442 528 1526 531
rect 1546 528 1686 531
rect 1710 528 1897 531
rect 1930 528 2062 531
rect 2098 528 2310 531
rect 2434 528 2497 531
rect 2570 528 2574 531
rect 2610 528 2630 531
rect 2634 528 2702 531
rect 2706 528 2726 531
rect 2806 528 2814 531
rect 2874 528 2910 531
rect 2954 528 3142 531
rect 3194 528 3222 531
rect 3378 528 3518 531
rect 3522 528 3534 531
rect 1710 522 1713 528
rect 66 518 110 521
rect 282 518 294 521
rect 370 518 390 521
rect 474 518 550 521
rect 618 518 622 521
rect 650 518 654 521
rect 770 518 806 521
rect 826 518 894 521
rect 930 518 934 521
rect 986 518 1270 521
rect 1274 518 1326 521
rect 1334 518 1417 521
rect 1426 518 1670 521
rect 1802 518 1862 521
rect 1874 518 1878 521
rect 1894 521 1897 528
rect 2494 522 2497 528
rect 2806 522 2809 528
rect 1894 518 1926 521
rect 1930 518 1950 521
rect 1982 518 1990 521
rect 1994 518 2054 521
rect 2522 518 2526 521
rect 2658 518 2662 521
rect 2674 518 2678 521
rect 2690 518 2702 521
rect 3098 518 3110 521
rect 3186 518 3198 521
rect 3202 518 3209 521
rect 3246 521 3249 528
rect 3218 518 3249 521
rect 258 508 350 511
rect 386 508 414 511
rect 458 508 614 511
rect 618 508 742 511
rect 810 508 814 511
rect 930 508 966 511
rect 1098 508 1182 511
rect 1202 508 1246 511
rect 1334 511 1337 518
rect 1322 508 1337 511
rect 1346 508 1358 511
rect 1362 508 1406 511
rect 1414 511 1417 518
rect 1414 508 1462 511
rect 1482 508 1590 511
rect 1618 508 1742 511
rect 1794 508 1974 511
rect 2202 508 2390 511
rect 2490 508 2590 511
rect 2594 508 2614 511
rect 2698 508 2702 511
rect 2778 508 2998 511
rect 3090 508 3198 511
rect 3530 508 3542 511
rect 992 503 994 507
rect 998 503 1001 507
rect 1006 503 1008 507
rect 1982 502 1985 508
rect 2024 503 2026 507
rect 2030 503 2033 507
rect 2038 503 2040 507
rect 3040 503 3042 507
rect 3046 503 3049 507
rect 3054 503 3056 507
rect 122 498 478 501
rect 482 498 558 501
rect 562 498 630 501
rect 642 498 726 501
rect 850 498 982 501
rect 1106 498 1206 501
rect 1274 498 1326 501
rect 1338 498 1430 501
rect 1442 498 1798 501
rect 1802 498 1822 501
rect 1898 498 1934 501
rect 2274 498 2382 501
rect 2514 498 2662 501
rect 2770 498 2774 501
rect 2818 498 2838 501
rect 3106 498 3150 501
rect 3154 498 3182 501
rect 3234 498 3278 501
rect 274 488 326 491
rect 478 488 486 491
rect 490 488 622 491
rect 654 488 662 491
rect 666 488 782 491
rect 862 488 870 491
rect 874 488 926 491
rect 1018 488 1054 491
rect 1090 488 1102 491
rect 1206 491 1209 498
rect 1206 488 1342 491
rect 1346 488 1406 491
rect 1434 488 1494 491
rect 1582 488 1590 491
rect 1594 488 1678 491
rect 1754 488 1822 491
rect 1834 488 1854 491
rect 1858 488 2014 491
rect 2018 488 2142 491
rect 2146 488 2401 491
rect 2562 488 2638 491
rect 2666 488 2710 491
rect 2742 488 2774 491
rect 2794 488 2814 491
rect 2830 488 3070 491
rect 3074 488 3094 491
rect 3202 488 3222 491
rect 3226 488 3390 491
rect 98 478 166 481
rect 262 481 265 488
rect 262 478 302 481
rect 338 478 406 481
rect 410 478 446 481
rect 474 478 614 481
rect 618 478 662 481
rect 682 478 686 481
rect 750 478 758 481
rect 762 478 870 481
rect 942 481 945 488
rect 922 478 945 481
rect 962 478 982 481
rect 986 478 1030 481
rect 1042 478 1150 481
rect 1162 478 1350 481
rect 1354 478 1542 481
rect 1550 481 1553 488
rect 2398 482 2401 488
rect 1550 478 1846 481
rect 1850 478 1870 481
rect 1874 478 1886 481
rect 2034 478 2046 481
rect 2066 478 2086 481
rect 2170 478 2174 481
rect 2258 478 2302 481
rect 2306 478 2318 481
rect 2330 478 2334 481
rect 2346 478 2350 481
rect 2402 478 2446 481
rect 2450 478 2566 481
rect 2642 478 2646 481
rect 2654 481 2657 488
rect 2654 478 2718 481
rect 2734 478 2737 488
rect 2742 482 2745 488
rect 2830 482 2833 488
rect 2770 478 2790 481
rect 2802 478 2806 481
rect 3034 478 3038 481
rect 3042 478 3217 481
rect 3226 478 3246 481
rect 3250 478 3334 481
rect 3410 478 3414 481
rect 26 468 30 471
rect 50 468 94 471
rect 206 471 209 478
rect 206 468 230 471
rect 282 468 286 471
rect 290 468 358 471
rect 362 468 390 471
rect 394 468 502 471
rect 506 468 510 471
rect 514 468 550 471
rect 554 468 582 471
rect 626 468 766 471
rect 770 468 822 471
rect 826 468 878 471
rect 938 468 942 471
rect 986 468 1078 471
rect 1106 468 1206 471
rect 1234 468 1326 471
rect 1394 468 1401 471
rect 1426 468 1510 471
rect 1530 468 1566 471
rect 1574 468 1582 471
rect 1586 468 1598 471
rect 1618 468 1646 471
rect 1834 468 1886 471
rect 1894 471 1897 478
rect 2182 472 2185 478
rect 1894 468 1990 471
rect 2010 468 2014 471
rect 2026 468 2110 471
rect 2138 468 2174 471
rect 2222 468 2246 471
rect 2306 468 2350 471
rect 2426 468 2430 471
rect 2602 468 2606 471
rect 2674 468 2814 471
rect 2938 468 3102 471
rect 3114 468 3118 471
rect 3146 468 3206 471
rect 3214 471 3217 478
rect 3214 468 3230 471
rect 3282 468 3310 471
rect 3314 468 3318 471
rect 3330 468 3334 471
rect 3338 468 3366 471
rect 3442 468 3534 471
rect 1398 462 1401 468
rect 26 458 286 461
rect 306 458 366 461
rect 370 458 374 461
rect 386 458 398 461
rect 410 458 414 461
rect 546 458 577 461
rect 602 458 622 461
rect 690 458 750 461
rect 786 458 854 461
rect 906 458 1062 461
rect 1146 458 1161 461
rect 1194 458 1257 461
rect 1290 458 1302 461
rect 1314 458 1342 461
rect 1482 458 1614 461
rect 1778 458 1782 461
rect 1866 458 1910 461
rect 1954 458 1966 461
rect 1994 458 2054 461
rect 2222 461 2225 468
rect 2074 458 2225 461
rect 2234 458 2294 461
rect 2322 458 2342 461
rect 2354 458 2390 461
rect 2458 458 2638 461
rect 2642 458 2846 461
rect 2962 458 2990 461
rect 3034 458 3089 461
rect 3114 458 3134 461
rect 3146 458 3326 461
rect 3330 458 3342 461
rect 3346 458 3374 461
rect 90 448 94 451
rect 170 448 558 451
rect 574 451 577 458
rect 870 452 873 458
rect 1094 452 1097 458
rect 1118 452 1121 458
rect 1158 452 1161 458
rect 1254 452 1257 458
rect 1414 452 1417 458
rect 574 448 630 451
rect 770 448 798 451
rect 858 448 862 451
rect 882 448 945 451
rect 710 442 713 448
rect 942 442 945 448
rect 950 448 990 451
rect 1010 448 1030 451
rect 1434 448 1513 451
rect 1522 448 1614 451
rect 1638 451 1641 458
rect 1638 448 1662 451
rect 1758 451 1761 458
rect 2310 452 2313 458
rect 1690 448 1761 451
rect 1794 448 1814 451
rect 1882 448 1902 451
rect 1974 448 2078 451
rect 2178 448 2238 451
rect 2250 448 2302 451
rect 2338 448 2502 451
rect 2538 448 2654 451
rect 2690 448 2694 451
rect 2746 448 2750 451
rect 2754 448 2798 451
rect 2882 448 2894 451
rect 2898 448 2902 451
rect 2910 451 2913 458
rect 2990 452 2993 458
rect 3086 452 3089 458
rect 2910 448 2926 451
rect 3114 448 3166 451
rect 3186 448 3278 451
rect 3306 448 3366 451
rect 3398 448 3470 451
rect 950 442 953 448
rect 178 438 182 441
rect 242 438 246 441
rect 314 438 342 441
rect 530 438 558 441
rect 610 438 646 441
rect 738 438 838 441
rect 1050 438 1054 441
rect 1090 438 1486 441
rect 1510 441 1513 448
rect 1510 438 1582 441
rect 1674 438 1742 441
rect 1786 438 1822 441
rect 1910 441 1913 448
rect 1850 438 1913 441
rect 1974 442 1977 448
rect 2078 441 2081 448
rect 2078 438 2150 441
rect 2166 441 2169 448
rect 2166 438 2318 441
rect 2370 438 2374 441
rect 2686 441 2689 448
rect 3398 442 3401 448
rect 2434 438 2689 441
rect 2722 438 2750 441
rect 2762 438 2790 441
rect 2794 438 2798 441
rect 2818 438 3030 441
rect 3074 438 3078 441
rect 3082 438 3241 441
rect 3266 438 3286 441
rect 206 432 209 438
rect 230 428 302 431
rect 306 428 430 431
rect 434 428 462 431
rect 518 431 521 438
rect 518 428 534 431
rect 586 428 686 431
rect 942 431 945 438
rect 942 428 1246 431
rect 1250 428 1294 431
rect 1410 428 1806 431
rect 1810 428 1870 431
rect 1922 428 2094 431
rect 2098 428 2166 431
rect 2170 428 2174 431
rect 2306 428 2454 431
rect 2594 428 2830 431
rect 2866 428 2886 431
rect 2890 428 2950 431
rect 3078 428 3086 431
rect 3090 428 3126 431
rect 3130 428 3134 431
rect 3146 428 3174 431
rect 3178 428 3182 431
rect 3238 431 3241 438
rect 3238 428 3334 431
rect 230 422 233 428
rect 30 418 230 421
rect 282 418 454 421
rect 530 418 574 421
rect 902 418 1070 421
rect 1074 418 1150 421
rect 1170 418 1174 421
rect 1434 418 1446 421
rect 1490 418 1550 421
rect 1626 418 1638 421
rect 1642 418 1654 421
rect 1698 418 1822 421
rect 1826 418 2022 421
rect 2058 418 2142 421
rect 2250 418 2390 421
rect 2394 418 2446 421
rect 2450 418 2502 421
rect 2626 418 2966 421
rect 2970 418 3062 421
rect 3066 418 3086 421
rect 3162 418 3190 421
rect 3194 418 3294 421
rect 3346 418 3422 421
rect 30 412 33 418
rect 226 408 230 411
rect 338 408 390 411
rect 514 408 614 411
rect 902 411 905 418
rect 714 408 905 411
rect 946 408 1326 411
rect 1394 408 1446 411
rect 1546 408 1926 411
rect 1930 408 1934 411
rect 1946 408 2118 411
rect 2142 411 2145 418
rect 2142 408 2246 411
rect 2330 408 2350 411
rect 2354 408 2366 411
rect 2794 408 2814 411
rect 2874 408 2902 411
rect 3002 408 3078 411
rect 3090 408 3406 411
rect 480 403 482 407
rect 486 403 489 407
rect 494 403 496 407
rect 1512 403 1514 407
rect 1518 403 1521 407
rect 1526 403 1528 407
rect 2536 403 2538 407
rect 2542 403 2545 407
rect 2550 403 2552 407
rect 370 398 462 401
rect 602 398 1022 401
rect 1130 398 1134 401
rect 1378 398 1478 401
rect 1634 398 1726 401
rect 1778 398 1878 401
rect 1922 398 2102 401
rect 2114 398 2230 401
rect 2282 398 2366 401
rect 2474 398 2478 401
rect 2578 398 2830 401
rect 2834 398 2942 401
rect 2954 398 3430 401
rect 242 388 414 391
rect 418 388 726 391
rect 730 388 790 391
rect 1066 388 1070 391
rect 1082 388 1134 391
rect 1210 388 1398 391
rect 1474 388 1718 391
rect 1722 388 1854 391
rect 1874 388 2950 391
rect 3002 388 3150 391
rect 3162 388 3182 391
rect 3242 388 3246 391
rect 3274 388 3302 391
rect 3330 388 3510 391
rect 2454 382 2457 388
rect 26 378 358 381
rect 450 378 766 381
rect 770 378 782 381
rect 786 378 854 381
rect 858 378 886 381
rect 890 378 1086 381
rect 1090 378 1198 381
rect 1202 378 1334 381
rect 1338 378 1542 381
rect 1546 378 1630 381
rect 1690 378 1878 381
rect 1898 378 1910 381
rect 1946 378 2006 381
rect 2010 378 2102 381
rect 2210 378 2358 381
rect 2478 378 3246 381
rect 3250 378 3286 381
rect 3442 378 3489 381
rect 586 368 590 371
rect 682 368 814 371
rect 882 368 902 371
rect 1018 368 1430 371
rect 1442 368 1446 371
rect 1514 368 1566 371
rect 1570 368 1670 371
rect 1678 371 1681 378
rect 2478 372 2481 378
rect 1678 368 1750 371
rect 1810 368 1902 371
rect 1906 368 1950 371
rect 1970 368 2478 371
rect 2610 368 2678 371
rect 2698 368 2814 371
rect 2826 368 2862 371
rect 3010 368 3030 371
rect 3042 368 3110 371
rect 3162 368 3190 371
rect 3406 371 3409 378
rect 3202 368 3409 371
rect 3486 372 3489 378
rect 638 362 641 368
rect 106 358 262 361
rect 266 358 270 361
rect 482 358 486 361
rect 554 358 582 361
rect 658 358 662 361
rect 870 361 873 368
rect 870 358 910 361
rect 930 358 934 361
rect 1038 358 1046 361
rect 1050 358 1070 361
rect 1182 358 1286 361
rect 1362 358 1406 361
rect 1450 358 1630 361
rect 1650 358 1790 361
rect 1946 358 1950 361
rect 1954 358 1982 361
rect 1994 358 2070 361
rect 2074 358 2182 361
rect 2210 358 2214 361
rect 2258 358 2278 361
rect 2282 358 2430 361
rect 2554 358 2614 361
rect 2682 358 2702 361
rect 2706 358 3078 361
rect 3082 358 3382 361
rect 3434 358 3510 361
rect -26 351 -22 352
rect 6 351 9 358
rect 614 352 617 358
rect -26 348 38 351
rect 42 348 62 351
rect 66 348 70 351
rect 138 348 174 351
rect 186 348 566 351
rect 578 348 582 351
rect 658 348 694 351
rect 698 348 702 351
rect 846 351 849 358
rect 1038 352 1041 358
rect 758 348 777 351
rect 846 348 910 351
rect 922 348 966 351
rect 970 348 998 351
rect 1026 348 1030 351
rect 1110 351 1113 358
rect 1182 352 1185 358
rect 1838 352 1841 358
rect 1058 348 1113 351
rect 1138 348 1142 351
rect 1154 348 1158 351
rect 1178 348 1182 351
rect 1210 348 1214 351
rect 1226 348 1230 351
rect 1258 348 1270 351
rect 1314 348 1350 351
rect 1394 348 1510 351
rect 1530 348 1542 351
rect 1618 348 1622 351
rect 1682 348 1694 351
rect 1738 348 1758 351
rect 1778 348 1782 351
rect 1810 348 1814 351
rect 1826 348 1830 351
rect 1846 351 1849 358
rect 1846 348 1862 351
rect 1898 348 1950 351
rect 1978 348 2022 351
rect 2106 348 2142 351
rect 2174 348 2198 351
rect 2206 348 2238 351
rect 2386 348 2430 351
rect 2442 348 2446 351
rect 2450 348 2574 351
rect 2586 348 2590 351
rect 2626 348 2654 351
rect 2686 348 2742 351
rect 2786 348 2806 351
rect 2842 348 2870 351
rect 2882 348 2886 351
rect 2962 348 3038 351
rect 3074 348 3078 351
rect 3098 348 3118 351
rect 3138 348 3158 351
rect 3194 348 3198 351
rect 3322 348 3342 351
rect 3374 348 3462 351
rect 3482 348 3542 351
rect 162 338 190 341
rect 246 338 278 341
rect 282 338 318 341
rect 322 338 334 341
rect 354 338 382 341
rect 506 338 526 341
rect 546 338 550 341
rect 566 341 569 348
rect 758 342 761 348
rect 774 342 777 348
rect 566 338 646 341
rect 650 338 710 341
rect 890 338 910 341
rect 922 338 934 341
rect 938 338 982 341
rect 1010 338 1174 341
rect 1178 338 1238 341
rect 1242 338 1262 341
rect 1466 338 1998 341
rect 2070 341 2073 348
rect 2174 342 2177 348
rect 2206 342 2209 348
rect 2686 342 2689 348
rect 2010 338 2102 341
rect 2130 338 2174 341
rect 2270 338 2302 341
rect 2402 338 2422 341
rect 2514 338 2534 341
rect 2578 338 2582 341
rect 2642 338 2686 341
rect 2722 338 2774 341
rect 2778 338 2822 341
rect 2878 341 2881 348
rect 2858 338 2881 341
rect 2898 338 2902 341
rect 2938 338 2942 341
rect 2978 338 2998 341
rect 3034 338 3102 341
rect 3122 338 3126 341
rect 3214 341 3217 348
rect 3374 342 3377 348
rect 3146 338 3217 341
rect 3234 338 3238 341
rect 3242 338 3350 341
rect 3402 338 3406 341
rect 3418 338 3510 341
rect 246 332 249 338
rect 186 328 206 331
rect 334 331 337 338
rect 870 332 873 338
rect 334 328 366 331
rect 378 328 454 331
rect 458 328 542 331
rect 570 328 622 331
rect 698 328 710 331
rect 746 328 774 331
rect 778 328 814 331
rect 970 328 998 331
rect 1374 331 1377 338
rect 2270 332 2273 338
rect 1002 328 1377 331
rect 1458 328 1462 331
rect 1498 328 1526 331
rect 1618 328 1702 331
rect 1802 328 1806 331
rect 1890 328 1910 331
rect 2026 328 2046 331
rect 2050 328 2078 331
rect 2114 328 2118 331
rect 2122 328 2190 331
rect 2266 328 2270 331
rect 2314 328 2326 331
rect 2330 328 2358 331
rect 2438 331 2441 338
rect 2418 328 2441 331
rect 2462 332 2465 338
rect 2498 328 2558 331
rect 2622 331 2625 338
rect 2622 328 2950 331
rect 2954 328 2958 331
rect 3074 328 3222 331
rect 3250 328 3262 331
rect 3290 328 3294 331
rect 3298 328 3318 331
rect 3426 328 3438 331
rect 178 318 182 321
rect 226 318 350 321
rect 394 318 398 321
rect 442 318 646 321
rect 650 318 678 321
rect 718 321 721 328
rect 1710 322 1713 328
rect 690 318 721 321
rect 746 318 750 321
rect 778 318 918 321
rect 946 318 1030 321
rect 1098 318 1118 321
rect 1202 318 1278 321
rect 1282 318 1382 321
rect 1426 318 1670 321
rect 1674 318 1686 321
rect 1794 318 2046 321
rect 2050 318 2222 321
rect 2226 318 2278 321
rect 2426 318 2486 321
rect 2578 318 2678 321
rect 2754 318 2790 321
rect 2810 318 2822 321
rect 2842 318 2974 321
rect 2990 321 2993 328
rect 2990 318 3038 321
rect 3058 318 3070 321
rect 3074 318 3102 321
rect 3186 318 3198 321
rect 3202 318 3254 321
rect 3266 318 3310 321
rect 3314 318 3358 321
rect 538 308 574 311
rect 586 308 598 311
rect 730 308 782 311
rect 802 308 838 311
rect 842 308 862 311
rect 1034 308 1246 311
rect 1258 308 1334 311
rect 1354 308 1366 311
rect 1370 308 1430 311
rect 1434 308 1470 311
rect 1482 308 1518 311
rect 1586 308 1662 311
rect 1666 308 1678 311
rect 1686 311 1689 318
rect 2574 312 2577 318
rect 1686 308 1726 311
rect 1818 308 1830 311
rect 1842 308 1862 311
rect 1866 308 1902 311
rect 1914 308 2006 311
rect 2162 308 2254 311
rect 2378 308 2470 311
rect 2714 308 2750 311
rect 2770 308 2774 311
rect 2898 308 2910 311
rect 2922 308 2958 311
rect 2978 308 2982 311
rect 3146 308 3166 311
rect 3170 308 3390 311
rect 992 303 994 307
rect 998 303 1001 307
rect 1006 303 1008 307
rect 2024 303 2026 307
rect 2030 303 2033 307
rect 2038 303 2040 307
rect 3040 303 3042 307
rect 3046 303 3049 307
rect 3054 303 3056 307
rect 282 298 294 301
rect 538 298 558 301
rect 826 298 830 301
rect 1114 298 1118 301
rect 1186 298 1254 301
rect 1338 298 1542 301
rect 1546 298 1854 301
rect 1906 298 1926 301
rect 1946 298 1998 301
rect 2002 298 2014 301
rect 2154 298 2166 301
rect 2346 298 2422 301
rect 2506 298 2542 301
rect 2562 298 2590 301
rect 2618 298 2630 301
rect 2714 298 2990 301
rect 3178 298 3270 301
rect 3362 298 3446 301
rect 3450 298 3470 301
rect 1326 292 1329 298
rect 206 288 214 291
rect 218 288 590 291
rect 594 288 670 291
rect 674 288 958 291
rect 962 288 1022 291
rect 1074 288 1094 291
rect 1194 288 1222 291
rect 1366 288 1374 291
rect 1378 288 1406 291
rect 1434 288 1702 291
rect 1706 288 1838 291
rect 1850 288 1854 291
rect 1866 288 2286 291
rect 2322 288 2358 291
rect 2366 288 2510 291
rect 2514 288 2518 291
rect 2738 288 2878 291
rect 2974 288 3006 291
rect 3250 288 3542 291
rect 86 281 89 288
rect 1110 282 1113 288
rect 1142 282 1145 288
rect 86 278 606 281
rect 666 278 806 281
rect 850 278 862 281
rect 930 278 934 281
rect 978 278 1038 281
rect 1130 278 1134 281
rect 1170 278 1182 281
rect 1274 278 1278 281
rect 1322 278 1366 281
rect 1458 278 1462 281
rect 1482 278 1550 281
rect 1586 278 1598 281
rect 1610 278 1614 281
rect 1626 278 1646 281
rect 1690 278 1694 281
rect 1706 278 1710 281
rect 1770 278 2094 281
rect 2098 278 2158 281
rect 2366 281 2369 288
rect 2298 278 2369 281
rect 2402 278 2430 281
rect 2562 278 2638 281
rect 2642 278 2710 281
rect 2918 281 2921 288
rect 2974 282 2977 288
rect 2826 278 2921 281
rect 2938 278 2950 281
rect 3130 278 3174 281
rect 3178 278 3238 281
rect 3338 278 3342 281
rect 170 268 214 271
rect 218 268 254 271
rect 314 268 358 271
rect 378 268 406 271
rect 410 268 462 271
rect 466 268 502 271
rect 618 268 622 271
rect 698 268 726 271
rect 746 268 750 271
rect 802 268 806 271
rect 1102 271 1105 278
rect 810 268 1286 271
rect 1290 268 1342 271
rect 1466 268 1470 271
rect 1490 268 1494 271
rect 1570 268 1574 271
rect 1586 268 1862 271
rect 1890 268 1910 271
rect 1914 268 1990 271
rect 2074 268 2094 271
rect 2138 268 2142 271
rect 2198 271 2201 278
rect 2806 272 2809 278
rect 3006 272 3009 278
rect 2194 268 2201 271
rect 2218 268 2302 271
rect 2314 268 2318 271
rect 2330 268 2334 271
rect 2386 268 2406 271
rect 2474 268 2486 271
rect 2490 268 2494 271
rect 2506 268 2510 271
rect 2522 268 2614 271
rect 2626 268 2630 271
rect 2674 268 2718 271
rect 2850 268 2902 271
rect 2906 268 2926 271
rect 3082 268 3142 271
rect 3146 268 3158 271
rect 3262 271 3265 278
rect 3166 268 3265 271
rect 3418 268 3430 271
rect 1542 262 1545 268
rect 66 258 662 261
rect 666 258 790 261
rect 810 258 814 261
rect 906 258 950 261
rect 1058 258 1150 261
rect 1178 258 1182 261
rect 1250 258 1262 261
rect 1306 258 1326 261
rect 1378 258 1409 261
rect 1426 258 1478 261
rect 1546 258 1598 261
rect 1610 258 1630 261
rect 1650 258 1718 261
rect 1746 258 1766 261
rect 1794 258 2022 261
rect 2066 258 2086 261
rect 2110 261 2113 268
rect 2110 258 2150 261
rect 2154 258 2222 261
rect 2226 258 2254 261
rect 2298 258 2382 261
rect 2394 258 2446 261
rect 2546 258 2657 261
rect 2666 258 2686 261
rect 2706 258 2726 261
rect 2730 258 2750 261
rect 2786 258 2806 261
rect 2818 258 2822 261
rect 2826 258 2854 261
rect 2874 258 2886 261
rect 2890 258 2934 261
rect 2998 261 3001 268
rect 3166 261 3169 268
rect 2998 258 3169 261
rect 3242 258 3318 261
rect 3426 258 3430 261
rect 3458 258 3486 261
rect 1406 252 1409 258
rect 1774 252 1777 258
rect 2478 252 2481 258
rect -26 251 -22 252
rect -26 248 6 251
rect 10 248 30 251
rect 34 248 70 251
rect 262 248 286 251
rect 322 248 526 251
rect 562 248 606 251
rect 610 248 614 251
rect 666 248 710 251
rect 754 248 758 251
rect 762 248 806 251
rect 810 248 990 251
rect 1042 248 1102 251
rect 1106 248 1110 251
rect 1122 248 1262 251
rect 1266 248 1270 251
rect 1290 248 1310 251
rect 1466 248 1558 251
rect 1570 248 1622 251
rect 1634 248 1646 251
rect 1670 248 1678 251
rect 1682 248 1758 251
rect 1802 248 1806 251
rect 1826 248 1830 251
rect 1874 248 1886 251
rect 1906 248 1926 251
rect 1930 248 2046 251
rect 2066 248 2086 251
rect 2098 248 2110 251
rect 2234 248 2238 251
rect 2242 248 2270 251
rect 2306 248 2398 251
rect 2402 248 2430 251
rect 2490 248 2566 251
rect 2570 248 2590 251
rect 2654 251 2657 258
rect 2654 248 2790 251
rect 2802 248 2950 251
rect 3066 248 3094 251
rect 3098 248 3126 251
rect 3170 248 3214 251
rect 3218 248 3278 251
rect 3482 248 3510 251
rect 3514 248 3558 251
rect 110 242 113 248
rect 262 242 265 248
rect 630 242 633 248
rect 638 242 641 248
rect 282 238 622 241
rect 642 238 726 241
rect 742 241 745 248
rect 742 238 758 241
rect 874 238 886 241
rect 938 238 1046 241
rect 1050 238 1094 241
rect 1098 238 1198 241
rect 1202 238 1238 241
rect 1286 241 1289 248
rect 1266 238 1289 241
rect 1322 238 1454 241
rect 1538 238 1550 241
rect 1610 238 1638 241
rect 1658 238 1846 241
rect 1850 238 1870 241
rect 1882 238 1910 241
rect 186 228 790 231
rect 850 228 902 231
rect 1130 228 1134 231
rect 1194 228 1286 231
rect 1290 228 1446 231
rect 1454 231 1457 238
rect 1454 228 1622 231
rect 1666 228 1790 231
rect 1850 228 1878 231
rect 1882 228 1918 231
rect 1958 231 1961 238
rect 1974 232 1977 238
rect 1982 232 1985 241
rect 1994 238 2206 241
rect 2286 241 2289 248
rect 2258 238 2289 241
rect 2378 238 2398 241
rect 2474 238 2558 241
rect 2594 238 2614 241
rect 2618 238 2678 241
rect 2682 238 2710 241
rect 2722 238 2942 241
rect 2946 238 3078 241
rect 3082 238 3150 241
rect 3402 238 3422 241
rect 3426 238 3494 241
rect 1958 228 1966 231
rect 1994 228 2030 231
rect 2130 228 2158 231
rect 2162 228 2318 231
rect 2338 228 2710 231
rect 2718 228 2862 231
rect 2866 228 2870 231
rect 2890 228 2902 231
rect 3026 228 3222 231
rect 2718 222 2721 228
rect 186 218 270 221
rect 274 218 318 221
rect 458 218 518 221
rect 522 218 838 221
rect 1194 218 1526 221
rect 1530 218 1582 221
rect 1682 218 2078 221
rect 2082 218 2286 221
rect 2290 218 2294 221
rect 2330 218 2510 221
rect 2530 218 2550 221
rect 2770 218 2774 221
rect 2994 218 3414 221
rect 926 212 929 218
rect 34 208 318 211
rect 586 208 614 211
rect 722 208 750 211
rect 754 208 822 211
rect 858 208 902 211
rect 930 208 1014 211
rect 1018 208 1022 211
rect 1186 208 1198 211
rect 1234 208 1246 211
rect 1258 208 1318 211
rect 1866 208 1934 211
rect 1946 208 2350 211
rect 2378 208 2382 211
rect 2394 208 2486 211
rect 2698 208 2958 211
rect 3194 208 3238 211
rect 3258 208 3542 211
rect 480 203 482 207
rect 486 203 489 207
rect 494 203 496 207
rect 1512 203 1514 207
rect 1518 203 1521 207
rect 1526 203 1528 207
rect 2536 203 2538 207
rect 2542 203 2545 207
rect 2550 203 2552 207
rect 154 198 446 201
rect 450 198 470 201
rect 506 198 566 201
rect 682 198 878 201
rect 938 198 998 201
rect 1034 198 1310 201
rect 1418 198 1430 201
rect 1730 198 1838 201
rect 1874 198 2270 201
rect 2282 198 2526 201
rect 2570 198 2737 201
rect 2746 198 2846 201
rect 2986 198 3470 201
rect 110 188 414 191
rect 418 188 542 191
rect 562 188 1206 191
rect 1210 188 2462 191
rect 2526 191 2529 198
rect 2526 188 2726 191
rect 2734 191 2737 198
rect 2734 188 2974 191
rect 2994 188 3022 191
rect 3050 188 3054 191
rect 3098 188 3382 191
rect 3390 188 3417 191
rect 110 182 113 188
rect 3390 182 3393 188
rect 3414 182 3417 188
rect 330 178 462 181
rect 466 178 470 181
rect 474 178 526 181
rect 530 178 590 181
rect 594 178 614 181
rect 618 178 774 181
rect 778 178 814 181
rect 818 178 838 181
rect 842 178 894 181
rect 914 178 1046 181
rect 1050 178 1118 181
rect 1122 178 1225 181
rect 1234 178 1350 181
rect 1450 178 1910 181
rect 1914 178 2166 181
rect 2178 178 2342 181
rect 2378 178 2382 181
rect 2610 178 2758 181
rect 2930 178 3230 181
rect 3274 178 3366 181
rect 54 171 57 178
rect 1222 172 1225 178
rect 54 168 190 171
rect 322 168 382 171
rect 386 168 430 171
rect 450 168 454 171
rect 462 168 574 171
rect 610 168 630 171
rect 638 168 758 171
rect 818 168 822 171
rect 834 168 870 171
rect 890 168 918 171
rect 938 168 1089 171
rect 1138 168 1142 171
rect 1178 168 1214 171
rect 1226 168 1406 171
rect 1410 168 1414 171
rect 1426 168 2862 171
rect 2866 168 2950 171
rect 2954 168 3110 171
rect 3154 168 3190 171
rect 3226 168 3294 171
rect 3394 168 3430 171
rect 298 158 302 161
rect 310 161 313 168
rect 310 158 334 161
rect 462 161 465 168
rect 338 158 465 161
rect 522 158 550 161
rect 638 161 641 168
rect 1086 162 1089 168
rect 554 158 641 161
rect 690 158 694 161
rect 706 158 710 161
rect 730 158 862 161
rect 882 158 886 161
rect 922 158 926 161
rect 954 158 958 161
rect 1090 158 1166 161
rect 1370 158 1542 161
rect 1562 158 1590 161
rect 1642 158 1678 161
rect 1914 158 1942 161
rect 2050 158 2054 161
rect 2058 158 2078 161
rect 2106 158 2126 161
rect 2186 158 2254 161
rect 2306 158 2350 161
rect 2442 158 2446 161
rect 2666 158 2670 161
rect 2682 158 2710 161
rect 2714 158 2734 161
rect 2842 158 2846 161
rect 2906 158 2910 161
rect 2922 158 2926 161
rect 2938 158 2942 161
rect 2954 158 2966 161
rect 2970 158 3062 161
rect 3170 158 3214 161
rect 3218 158 3246 161
rect 3306 158 3318 161
rect 3402 158 3550 161
rect 1334 152 1337 158
rect 1342 152 1345 158
rect 34 148 542 151
rect 546 148 582 151
rect 586 148 1246 151
rect 1250 148 1302 151
rect 1354 148 1358 151
rect 1362 148 1414 151
rect 1422 148 1446 151
rect 1490 148 1534 151
rect 1546 148 1670 151
rect 1674 148 1694 151
rect 1742 151 1745 158
rect 2142 152 2145 158
rect 1706 148 1745 151
rect 1762 148 1806 151
rect 1874 148 1950 151
rect 1954 148 2006 151
rect 2050 148 2110 151
rect 2170 148 2190 151
rect 2210 148 2294 151
rect 2330 148 2350 151
rect 2362 148 2366 151
rect 2418 148 2422 151
rect 2506 148 2654 151
rect 2678 148 2790 151
rect 2794 148 2806 151
rect 2826 148 2830 151
rect 2870 151 2873 158
rect 2858 148 2873 151
rect 2882 148 2886 151
rect 2898 148 3038 151
rect 3042 148 3046 151
rect 3098 148 3102 151
rect 3142 151 3145 158
rect 3114 148 3145 151
rect 3178 148 3182 151
rect 3186 148 3278 151
rect 3290 148 3342 151
rect 3386 148 3406 151
rect 106 138 118 141
rect 138 138 166 141
rect 170 138 198 141
rect 218 138 278 141
rect 362 138 502 141
rect 506 138 510 141
rect 522 138 574 141
rect 626 138 638 141
rect 658 138 662 141
rect 722 138 726 141
rect 738 138 742 141
rect 770 138 774 141
rect 810 138 838 141
rect 866 138 950 141
rect 966 138 1054 141
rect 1114 138 1118 141
rect 1162 138 1166 141
rect 1186 138 1190 141
rect 1218 138 1230 141
rect 1266 138 1270 141
rect 1290 138 1342 141
rect 1382 138 1390 141
rect 1422 141 1425 148
rect 1394 138 1425 141
rect 1434 138 1438 141
rect 1458 138 1494 141
rect 1562 138 1590 141
rect 1602 138 1654 141
rect 1666 138 1798 141
rect 1814 141 1817 148
rect 1814 138 1862 141
rect 1866 138 1910 141
rect 1970 138 2078 141
rect 2122 138 2158 141
rect 2162 138 2206 141
rect 2210 138 2230 141
rect 2274 138 2406 141
rect 2426 138 2438 141
rect 2678 141 2681 148
rect 2514 138 2681 141
rect 2770 138 2774 141
rect 2778 138 2886 141
rect 2890 138 2902 141
rect 2946 138 2982 141
rect 3098 138 3182 141
rect 3186 138 3342 141
rect 3346 138 3358 141
rect 3370 138 3382 141
rect 3386 138 3478 141
rect 214 132 217 138
rect 966 132 969 138
rect 290 128 430 131
rect 434 128 577 131
rect 586 128 702 131
rect 722 128 734 131
rect 762 128 926 131
rect 930 128 966 131
rect 986 128 1078 131
rect 1082 128 1177 131
rect 1234 128 1358 131
rect 1374 131 1377 138
rect 1374 128 1390 131
rect 1458 128 1526 131
rect 1562 128 1582 131
rect 1586 128 1590 131
rect 1706 128 1710 131
rect 1770 128 1854 131
rect 1858 128 1886 131
rect 1938 128 2062 131
rect 2074 128 2110 131
rect 2114 128 2126 131
rect 2134 128 2142 131
rect 2154 128 2166 131
rect 2182 128 2398 131
rect 2410 128 2422 131
rect 2486 131 2489 138
rect 2750 132 2753 138
rect 3022 132 3025 138
rect 3518 132 3521 138
rect 2482 128 2489 131
rect 2498 128 2502 131
rect 2594 128 2646 131
rect 2650 128 2694 131
rect 2810 128 2814 131
rect 2822 128 2830 131
rect 2834 128 2870 131
rect 3074 128 3110 131
rect 3122 128 3286 131
rect 3298 128 3310 131
rect 3322 128 3326 131
rect 3346 128 3350 131
rect 3362 128 3366 131
rect 3426 128 3454 131
rect 378 118 382 121
rect 442 118 446 121
rect 574 121 577 128
rect 1174 122 1177 128
rect 2182 122 2185 128
rect 250 108 366 111
rect 438 111 441 118
rect 378 108 441 111
rect 454 112 457 121
rect 574 118 582 121
rect 586 118 670 121
rect 674 118 766 121
rect 810 118 894 121
rect 898 118 1150 121
rect 1178 118 1190 121
rect 1242 118 1262 121
rect 1266 118 1302 121
rect 1322 118 1382 121
rect 1402 118 1486 121
rect 1490 118 1550 121
rect 1554 118 1614 121
rect 1730 118 1798 121
rect 1810 118 1926 121
rect 1978 118 2006 121
rect 2010 118 2110 121
rect 2114 118 2174 121
rect 2242 118 2478 121
rect 2490 118 2566 121
rect 2570 118 2622 121
rect 2658 118 2766 121
rect 2794 118 2886 121
rect 2970 118 3134 121
rect 3138 118 3158 121
rect 3226 118 3302 121
rect 3314 118 3486 121
rect 3490 118 3526 121
rect 514 108 558 111
rect 626 108 630 111
rect 794 108 822 111
rect 874 108 878 111
rect 914 108 950 111
rect 1018 108 1110 111
rect 1114 108 1310 111
rect 1314 108 1766 111
rect 1786 108 1814 111
rect 1834 108 1942 111
rect 2098 108 2166 111
rect 2194 108 2246 111
rect 2258 108 2318 111
rect 2330 108 2334 111
rect 2354 108 2358 111
rect 2378 108 2662 111
rect 2778 108 2886 111
rect 2898 108 3014 111
rect 3154 108 3174 111
rect 3178 108 3334 111
rect 3378 108 3454 111
rect 982 102 985 108
rect 992 103 994 107
rect 998 103 1001 107
rect 1006 103 1008 107
rect 2024 103 2026 107
rect 2030 103 2033 107
rect 2038 103 2040 107
rect 3040 103 3042 107
rect 3046 103 3049 107
rect 3054 103 3056 107
rect 266 98 270 101
rect 282 98 542 101
rect 626 98 638 101
rect 826 98 862 101
rect 866 98 886 101
rect 946 98 974 101
rect 1026 98 1062 101
rect 1066 98 1102 101
rect 1162 98 1382 101
rect 1386 98 1534 101
rect 1538 98 1638 101
rect 1642 98 1670 101
rect 1674 98 1734 101
rect 1770 98 1798 101
rect 1818 98 1942 101
rect 1946 98 1974 101
rect 2050 98 2118 101
rect 2282 98 2286 101
rect 2298 98 2326 101
rect 2402 98 2406 101
rect 2418 98 2446 101
rect 2458 98 2606 101
rect 2618 98 2670 101
rect 2682 98 2958 101
rect 3010 98 3030 101
rect 3066 98 3094 101
rect 3106 98 3310 101
rect 3322 98 3326 101
rect 3346 98 3430 101
rect 3454 98 3462 101
rect 3466 98 3510 101
rect 150 88 158 91
rect 162 88 246 91
rect 250 88 342 91
rect 394 88 398 91
rect 434 88 550 91
rect 554 88 558 91
rect 570 88 606 91
rect 698 88 718 91
rect 730 88 734 91
rect 750 88 758 91
rect 762 88 782 91
rect 794 88 1126 91
rect 1130 88 1198 91
rect 1250 88 2126 91
rect 2130 88 2502 91
rect 2506 88 2566 91
rect 2586 88 2590 91
rect 2630 88 2710 91
rect 2722 88 2758 91
rect 2762 88 3014 91
rect 3018 88 3134 91
rect 3454 91 3457 98
rect 3194 88 3457 91
rect 54 81 57 88
rect 54 78 102 81
rect 118 81 121 88
rect 2630 82 2633 88
rect 3462 82 3465 88
rect 118 78 510 81
rect 514 78 937 81
rect 946 78 990 81
rect 1026 78 1038 81
rect 1058 78 1070 81
rect 1074 78 1182 81
rect 1210 78 1214 81
rect 1290 78 1294 81
rect 1362 78 1398 81
rect 1418 78 1446 81
rect 1466 78 1489 81
rect 1506 78 1558 81
rect 1618 78 1686 81
rect 1698 78 1846 81
rect 1850 78 1870 81
rect 1882 78 1886 81
rect 1898 78 1902 81
rect 1922 78 1926 81
rect 1962 78 1966 81
rect 1986 78 1990 81
rect 2010 78 2014 81
rect 2034 78 2046 81
rect 2058 78 2062 81
rect 2194 78 2438 81
rect 2466 78 2478 81
rect 2486 78 2614 81
rect 2690 78 2694 81
rect 2802 78 2806 81
rect 2890 78 2918 81
rect 2942 78 2977 81
rect 34 68 422 71
rect 442 68 478 71
rect 546 68 614 71
rect 618 68 670 71
rect 674 68 806 71
rect 834 68 838 71
rect 866 68 870 71
rect 934 71 937 78
rect 934 68 958 71
rect 962 68 966 71
rect 970 68 1078 71
rect 1090 68 1094 71
rect 1146 68 1182 71
rect 1186 68 1206 71
rect 1226 68 1238 71
rect 1290 68 1294 71
rect 1350 71 1353 78
rect 1486 72 1489 78
rect 1314 68 1430 71
rect 1434 68 1470 71
rect 1474 68 1478 71
rect 1498 68 1518 71
rect 1522 68 2158 71
rect 2210 68 2230 71
rect 2290 68 2318 71
rect 2486 71 2489 78
rect 2750 72 2753 78
rect 2862 72 2865 78
rect 2942 72 2945 78
rect 2974 72 2977 78
rect 3050 78 3206 81
rect 3290 78 3294 81
rect 3346 78 3438 81
rect 3030 72 3033 78
rect 3038 72 3041 78
rect 3478 72 3481 78
rect 2322 68 2489 71
rect 2562 68 2590 71
rect 2594 68 2646 71
rect 2682 68 2726 71
rect 2810 68 2854 71
rect 2930 68 2934 71
rect 2954 68 2966 71
rect 3138 68 3150 71
rect 3154 68 3206 71
rect 3210 68 3310 71
rect 3322 68 3326 71
rect 3338 68 3342 71
rect 2262 62 2265 68
rect 10 58 46 61
rect 74 58 206 61
rect 234 58 686 61
rect 690 58 822 61
rect 826 58 998 61
rect 1034 58 1094 61
rect 1098 58 1102 61
rect 1218 58 1222 61
rect 1250 58 1278 61
rect 1322 58 1342 61
rect 1354 58 1358 61
rect 1370 58 1374 61
rect 1426 58 1430 61
rect 1442 58 1446 61
rect 1450 58 1478 61
rect 1506 58 1526 61
rect 1530 58 1614 61
rect 1690 58 1742 61
rect 1746 58 1822 61
rect 1826 58 1998 61
rect 2010 58 2118 61
rect 2146 58 2198 61
rect 2218 58 2222 61
rect 2234 58 2238 61
rect 2242 58 2254 61
rect 2266 58 2326 61
rect 2330 58 2334 61
rect 2362 58 2366 61
rect 2386 58 2390 61
rect 2442 58 2454 61
rect 2466 58 2542 61
rect 2674 58 2702 61
rect 2722 58 2734 61
rect 2738 58 2774 61
rect 2786 58 3374 61
rect 3538 58 3550 61
rect 74 48 102 51
rect 106 48 222 51
rect 226 48 246 51
rect 262 48 350 51
rect 370 48 478 51
rect 482 48 486 51
rect 562 48 566 51
rect 610 48 654 51
rect 666 48 670 51
rect 674 48 766 51
rect 770 48 798 51
rect 850 48 854 51
rect 874 48 1022 51
rect 1118 51 1121 58
rect 1030 48 1222 51
rect 1234 48 1238 51
rect 1250 48 1406 51
rect 1442 48 1454 51
rect 1482 48 1622 51
rect 1630 51 1633 58
rect 1626 48 1633 51
rect 1642 48 1782 51
rect 1810 48 1814 51
rect 1842 48 1902 51
rect 1906 48 1910 51
rect 1914 48 1950 51
rect 2118 51 2121 58
rect 2462 52 2465 58
rect 2118 48 2334 51
rect 2338 48 2374 51
rect 2378 48 2406 51
rect 2410 48 2430 51
rect 2554 48 2582 51
rect 2602 48 2614 51
rect 2842 48 2966 51
rect 2978 48 3046 51
rect 3138 48 3142 51
rect 3234 48 3398 51
rect 3590 48 3594 52
rect 262 42 265 48
rect 86 38 230 41
rect 314 38 390 41
rect 394 38 726 41
rect 786 38 790 41
rect 818 38 878 41
rect 1030 41 1033 48
rect 882 38 1033 41
rect 1042 38 1086 41
rect 1162 38 1566 41
rect 1570 38 1702 41
rect 1706 38 1774 41
rect 1778 38 1830 41
rect 1838 38 1846 41
rect 1850 38 1870 41
rect 1874 38 1990 41
rect 1994 38 2294 41
rect 2306 38 2590 41
rect 2866 38 2886 41
rect 2954 38 2958 41
rect 86 32 89 38
rect 410 28 438 31
rect 442 28 449 31
rect 458 28 558 31
rect 698 28 702 31
rect 714 28 726 31
rect 786 28 1062 31
rect 1066 28 1102 31
rect 2302 31 2305 38
rect 1106 28 2305 31
rect 2362 28 2574 31
rect 2606 31 2609 38
rect 2966 32 2969 41
rect 2978 38 3078 41
rect 3082 38 3158 41
rect 3218 38 3254 41
rect 3590 41 3593 48
rect 3310 38 3593 41
rect 3310 32 3313 38
rect 2606 28 2918 31
rect 602 18 606 21
rect 650 18 654 21
rect 666 18 694 21
rect 698 18 1158 21
rect 1558 18 1566 21
rect 1570 18 1646 21
rect 2210 18 2422 21
rect 2570 18 2582 21
rect 2682 18 2686 21
rect 2858 18 2982 21
rect 2986 18 2990 21
rect 2994 18 3006 21
rect 1214 12 1217 18
rect 1486 12 1489 18
rect 2766 12 2769 18
rect 274 8 286 11
rect 538 8 622 11
rect 626 8 726 11
rect 810 8 814 11
rect 890 8 974 11
rect 1050 8 1054 11
rect 1266 8 1270 11
rect 1546 8 1550 11
rect 1602 8 1614 11
rect 2338 8 2342 11
rect 2370 8 2374 11
rect 2418 8 2422 11
rect 2706 8 2758 11
rect 2850 8 2862 11
rect 2914 8 3078 11
rect 3338 8 3350 11
rect 480 3 482 7
rect 486 3 489 7
rect 494 3 496 7
rect 1512 3 1514 7
rect 1518 3 1521 7
rect 1526 3 1528 7
rect 2536 3 2538 7
rect 2542 3 2545 7
rect 2550 3 2552 7
<< m4contact >>
rect 994 3303 998 3307
rect 1002 3303 1005 3307
rect 1005 3303 1006 3307
rect 2026 3303 2030 3307
rect 2034 3303 2037 3307
rect 2037 3303 2038 3307
rect 3042 3303 3046 3307
rect 3050 3303 3053 3307
rect 3053 3303 3054 3307
rect 686 3298 690 3302
rect 1134 3298 1138 3302
rect 1294 3298 1298 3302
rect 1374 3298 1378 3302
rect 1406 3298 1410 3302
rect 1542 3298 1546 3302
rect 1654 3298 1658 3302
rect 1718 3298 1722 3302
rect 1734 3298 1738 3302
rect 1918 3298 1922 3302
rect 1998 3298 2002 3302
rect 2198 3298 2202 3302
rect 2254 3298 2258 3302
rect 2462 3298 2466 3302
rect 2518 3298 2522 3302
rect 2638 3298 2642 3302
rect 2646 3298 2650 3302
rect 2806 3298 2810 3302
rect 3078 3298 3082 3302
rect 606 3288 610 3292
rect 670 3288 674 3292
rect 1022 3288 1026 3292
rect 1054 3288 1058 3292
rect 1230 3288 1234 3292
rect 1598 3288 1602 3292
rect 2158 3288 2162 3292
rect 2174 3288 2178 3292
rect 2230 3288 2234 3292
rect 2246 3288 2250 3292
rect 2790 3288 2794 3292
rect 2926 3288 2930 3292
rect 630 3278 634 3282
rect 886 3278 890 3282
rect 1534 3278 1538 3282
rect 3510 3278 3514 3282
rect 718 3268 722 3272
rect 1454 3268 1458 3272
rect 1646 3268 1650 3272
rect 1702 3268 1706 3272
rect 2574 3268 2578 3272
rect 2854 3268 2858 3272
rect 3294 3268 3298 3272
rect 3310 3268 3314 3272
rect 3390 3268 3394 3272
rect 3438 3268 3442 3272
rect 3518 3268 3522 3272
rect 1286 3258 1290 3262
rect 1534 3258 1538 3262
rect 1838 3258 1842 3262
rect 2038 3258 2042 3262
rect 2214 3258 2218 3262
rect 2310 3258 2314 3262
rect 2470 3258 2474 3262
rect 2678 3258 2682 3262
rect 2758 3258 2762 3262
rect 2918 3258 2922 3262
rect 3094 3258 3098 3262
rect 3126 3258 3130 3262
rect 3174 3258 3178 3262
rect 3366 3258 3370 3262
rect 3374 3258 3378 3262
rect 3398 3258 3402 3262
rect 3454 3258 3458 3262
rect 614 3248 618 3252
rect 1078 3248 1082 3252
rect 1246 3248 1250 3252
rect 1422 3248 1426 3252
rect 2502 3248 2506 3252
rect 3446 3248 3450 3252
rect 3550 3248 3554 3252
rect 1286 3238 1290 3242
rect 734 3228 738 3232
rect 1430 3228 1434 3232
rect 3502 3228 3506 3232
rect 1078 3218 1082 3222
rect 1950 3218 1954 3222
rect 1878 3208 1882 3212
rect 2454 3208 2458 3212
rect 482 3203 486 3207
rect 490 3203 493 3207
rect 493 3203 494 3207
rect 1514 3203 1518 3207
rect 1522 3203 1525 3207
rect 1525 3203 1526 3207
rect 2538 3203 2542 3207
rect 2546 3203 2549 3207
rect 2549 3203 2550 3207
rect 1502 3198 1506 3202
rect 1670 3198 1674 3202
rect 1958 3198 1962 3202
rect 3358 3198 3362 3202
rect 3214 3188 3218 3192
rect 3102 3178 3106 3182
rect 758 3168 762 3172
rect 838 3168 842 3172
rect 1742 3168 1746 3172
rect 1198 3158 1202 3162
rect 1286 3158 1290 3162
rect 2486 3158 2490 3162
rect 2710 3158 2714 3162
rect 3294 3158 3298 3162
rect 310 3148 314 3152
rect 854 3148 858 3152
rect 902 3148 906 3152
rect 1142 3148 1146 3152
rect 1350 3148 1354 3152
rect 1462 3148 1466 3152
rect 1862 3148 1866 3152
rect 1910 3148 1914 3152
rect 2062 3148 2066 3152
rect 2782 3148 2786 3152
rect 3326 3148 3330 3152
rect 974 3138 978 3142
rect 1134 3138 1138 3142
rect 1342 3138 1346 3142
rect 1646 3138 1650 3142
rect 2190 3138 2194 3142
rect 2310 3138 2314 3142
rect 2678 3138 2682 3142
rect 2774 3138 2778 3142
rect 2998 3138 3002 3142
rect 3470 3138 3474 3142
rect 3494 3138 3498 3142
rect 206 3128 210 3132
rect 1398 3128 1402 3132
rect 1446 3128 1450 3132
rect 1662 3128 1666 3132
rect 2174 3128 2178 3132
rect 2262 3128 2266 3132
rect 2470 3128 2474 3132
rect 1014 3118 1018 3122
rect 1030 3118 1034 3122
rect 1102 3118 1106 3122
rect 1110 3118 1114 3122
rect 1990 3118 1994 3122
rect 2222 3118 2226 3122
rect 2526 3118 2530 3122
rect 710 3108 714 3112
rect 798 3108 802 3112
rect 918 3108 922 3112
rect 1374 3108 1378 3112
rect 1814 3108 1818 3112
rect 1966 3108 1970 3112
rect 2206 3108 2210 3112
rect 2214 3108 2218 3112
rect 2366 3108 2370 3112
rect 3174 3108 3178 3112
rect 3302 3108 3306 3112
rect 994 3103 998 3107
rect 1002 3103 1005 3107
rect 1005 3103 1006 3107
rect 2026 3103 2030 3107
rect 2034 3103 2037 3107
rect 2037 3103 2038 3107
rect 3042 3103 3046 3107
rect 3050 3103 3053 3107
rect 3053 3103 3054 3107
rect 1014 3098 1018 3102
rect 614 3088 618 3092
rect 1622 3088 1626 3092
rect 1862 3088 1866 3092
rect 2014 3088 2018 3092
rect 2214 3088 2218 3092
rect 2318 3088 2322 3092
rect 606 3078 610 3082
rect 902 3078 906 3082
rect 1126 3078 1130 3082
rect 1150 3078 1154 3082
rect 1214 3078 1218 3082
rect 1294 3078 1298 3082
rect 2086 3078 2090 3082
rect 2166 3078 2170 3082
rect 2222 3078 2226 3082
rect 2438 3078 2442 3082
rect 2854 3078 2858 3082
rect 166 3068 170 3072
rect 1622 3068 1626 3072
rect 1750 3068 1754 3072
rect 1830 3068 1834 3072
rect 2094 3068 2098 3072
rect 2174 3068 2178 3072
rect 2510 3068 2514 3072
rect 334 3058 338 3062
rect 566 3058 570 3062
rect 854 3058 858 3062
rect 1334 3058 1338 3062
rect 1782 3058 1786 3062
rect 2062 3058 2066 3062
rect 2182 3058 2186 3062
rect 2350 3058 2354 3062
rect 2510 3058 2514 3062
rect 2782 3058 2786 3062
rect 2910 3058 2914 3062
rect 342 3048 346 3052
rect 590 3048 594 3052
rect 942 3048 946 3052
rect 1470 3048 1474 3052
rect 1494 3048 1498 3052
rect 1902 3048 1906 3052
rect 1990 3048 1994 3052
rect 2126 3048 2130 3052
rect 2590 3048 2594 3052
rect 3086 3048 3090 3052
rect 382 3038 386 3042
rect 598 3038 602 3042
rect 1134 3038 1138 3042
rect 1318 3038 1322 3042
rect 2190 3038 2194 3042
rect 2318 3038 2322 3042
rect 2766 3038 2770 3042
rect 542 3028 546 3032
rect 694 3028 698 3032
rect 726 3028 730 3032
rect 830 3028 834 3032
rect 1702 3028 1706 3032
rect 2446 3028 2450 3032
rect 718 3018 722 3022
rect 1230 3018 1234 3022
rect 2270 3018 2274 3022
rect 1150 3008 1154 3012
rect 2558 3008 2562 3012
rect 3310 3008 3314 3012
rect 482 3003 486 3007
rect 490 3003 493 3007
rect 493 3003 494 3007
rect 1514 3003 1518 3007
rect 1522 3003 1525 3007
rect 1525 3003 1526 3007
rect 2538 3003 2542 3007
rect 2546 3003 2549 3007
rect 2549 3003 2550 3007
rect 758 2998 762 3002
rect 1102 2998 1106 3002
rect 1478 2998 1482 3002
rect 1502 2998 1506 3002
rect 2470 2998 2474 3002
rect 2990 2998 2994 3002
rect 854 2988 858 2992
rect 1054 2988 1058 2992
rect 1246 2988 1250 2992
rect 1590 2988 1594 2992
rect 2238 2988 2242 2992
rect 3006 2988 3010 2992
rect 654 2978 658 2982
rect 886 2978 890 2982
rect 926 2978 930 2982
rect 1358 2978 1362 2982
rect 1462 2978 1466 2982
rect 2246 2978 2250 2982
rect 3510 2978 3514 2982
rect 110 2968 114 2972
rect 1118 2968 1122 2972
rect 1230 2968 1234 2972
rect 1438 2958 1442 2962
rect 1734 2958 1738 2962
rect 3206 2958 3210 2962
rect 3270 2958 3274 2962
rect 3542 2958 3546 2962
rect 230 2948 234 2952
rect 262 2948 266 2952
rect 670 2948 674 2952
rect 734 2948 738 2952
rect 846 2948 850 2952
rect 1014 2948 1018 2952
rect 1046 2948 1050 2952
rect 1062 2948 1066 2952
rect 1094 2948 1098 2952
rect 2046 2948 2050 2952
rect 2174 2948 2178 2952
rect 2198 2948 2202 2952
rect 2366 2948 2370 2952
rect 2526 2948 2530 2952
rect 126 2938 130 2942
rect 742 2938 746 2942
rect 814 2938 818 2942
rect 998 2938 1002 2942
rect 1126 2938 1130 2942
rect 1230 2938 1234 2942
rect 430 2928 434 2932
rect 630 2928 634 2932
rect 766 2928 770 2932
rect 774 2928 778 2932
rect 798 2928 802 2932
rect 830 2928 834 2932
rect 862 2928 866 2932
rect 918 2928 922 2932
rect 966 2928 970 2932
rect 974 2928 978 2932
rect 1006 2928 1010 2932
rect 1766 2938 1770 2942
rect 1822 2938 1826 2942
rect 2030 2938 2034 2942
rect 2502 2938 2506 2942
rect 2878 2938 2882 2942
rect 3422 2938 3426 2942
rect 1182 2928 1186 2932
rect 1358 2928 1362 2932
rect 1438 2928 1442 2932
rect 1646 2928 1650 2932
rect 1798 2928 1802 2932
rect 1862 2928 1866 2932
rect 1878 2928 1882 2932
rect 1934 2928 1938 2932
rect 2014 2928 2018 2932
rect 2078 2928 2082 2932
rect 2502 2928 2506 2932
rect 2934 2928 2938 2932
rect 3270 2928 3274 2932
rect 46 2918 50 2922
rect 1318 2918 1322 2922
rect 1350 2918 1354 2922
rect 1382 2918 1386 2922
rect 1606 2918 1610 2922
rect 1622 2918 1626 2922
rect 1734 2918 1738 2922
rect 3118 2918 3122 2922
rect 134 2908 138 2912
rect 1038 2908 1042 2912
rect 1262 2908 1266 2912
rect 1910 2908 1914 2912
rect 2118 2908 2122 2912
rect 994 2903 998 2907
rect 1002 2903 1005 2907
rect 1005 2903 1006 2907
rect 414 2898 418 2902
rect 446 2898 450 2902
rect 966 2898 970 2902
rect 1086 2898 1090 2902
rect 1110 2898 1114 2902
rect 1470 2898 1474 2902
rect 2026 2903 2030 2907
rect 2034 2903 2037 2907
rect 2037 2903 2038 2907
rect 3042 2903 3046 2907
rect 3050 2903 3053 2907
rect 3053 2903 3054 2907
rect 1814 2898 1818 2902
rect 1926 2898 1930 2902
rect 1982 2898 1986 2902
rect 2470 2898 2474 2902
rect 2774 2898 2778 2902
rect 3518 2898 3522 2902
rect 3534 2898 3538 2902
rect 286 2888 290 2892
rect 630 2888 634 2892
rect 726 2888 730 2892
rect 1054 2888 1058 2892
rect 1078 2888 1082 2892
rect 1118 2888 1122 2892
rect 1142 2888 1146 2892
rect 1262 2888 1266 2892
rect 1302 2888 1306 2892
rect 3198 2888 3202 2892
rect 3446 2888 3450 2892
rect 238 2878 242 2882
rect 278 2878 282 2882
rect 398 2878 402 2882
rect 558 2878 562 2882
rect 662 2878 666 2882
rect 734 2878 738 2882
rect 1062 2878 1066 2882
rect 1286 2878 1290 2882
rect 1478 2878 1482 2882
rect 1550 2878 1554 2882
rect 1662 2878 1666 2882
rect 1846 2878 1850 2882
rect 1886 2878 1890 2882
rect 2110 2878 2114 2882
rect 2358 2878 2362 2882
rect 2454 2878 2458 2882
rect 2606 2878 2610 2882
rect 3318 2878 3322 2882
rect 3342 2878 3346 2882
rect 3486 2878 3490 2882
rect 366 2868 370 2872
rect 422 2868 426 2872
rect 734 2868 738 2872
rect 758 2868 762 2872
rect 886 2868 890 2872
rect 902 2868 906 2872
rect 934 2868 938 2872
rect 1134 2868 1138 2872
rect 1374 2868 1378 2872
rect 1622 2868 1626 2872
rect 1726 2868 1730 2872
rect 2150 2868 2154 2872
rect 2254 2868 2258 2872
rect 2478 2868 2482 2872
rect 2494 2868 2498 2872
rect 2598 2868 2602 2872
rect 2790 2868 2794 2872
rect 2998 2868 3002 2872
rect 3366 2868 3370 2872
rect 3526 2868 3530 2872
rect 30 2858 34 2862
rect 126 2858 130 2862
rect 510 2858 514 2862
rect 638 2858 642 2862
rect 854 2858 858 2862
rect 1126 2858 1130 2862
rect 1382 2858 1386 2862
rect 1486 2858 1490 2862
rect 1838 2858 1842 2862
rect 1902 2858 1906 2862
rect 1918 2858 1922 2862
rect 1998 2858 2002 2862
rect 2078 2858 2082 2862
rect 2214 2858 2218 2862
rect 2286 2858 2290 2862
rect 2566 2858 2570 2862
rect 2998 2858 3002 2862
rect 294 2848 298 2852
rect 310 2848 314 2852
rect 358 2848 362 2852
rect 1326 2848 1330 2852
rect 1654 2848 1658 2852
rect 1694 2848 1698 2852
rect 1774 2848 1778 2852
rect 1790 2848 1794 2852
rect 1942 2848 1946 2852
rect 1958 2848 1962 2852
rect 2574 2848 2578 2852
rect 2806 2848 2810 2852
rect 3262 2848 3266 2852
rect 3350 2848 3354 2852
rect 46 2838 50 2842
rect 1414 2838 1418 2842
rect 1590 2838 1594 2842
rect 2494 2838 2498 2842
rect 2742 2838 2746 2842
rect 3134 2838 3138 2842
rect 3334 2838 3338 2842
rect 278 2828 282 2832
rect 430 2828 434 2832
rect 526 2828 530 2832
rect 1070 2828 1074 2832
rect 1830 2828 1834 2832
rect 2182 2828 2186 2832
rect 2206 2828 2210 2832
rect 2806 2828 2810 2832
rect 102 2818 106 2822
rect 1246 2818 1250 2822
rect 1966 2818 1970 2822
rect 2158 2818 2162 2822
rect 2478 2818 2482 2822
rect 2486 2818 2490 2822
rect 3318 2818 3322 2822
rect 662 2808 666 2812
rect 966 2808 970 2812
rect 1318 2808 1322 2812
rect 1350 2808 1354 2812
rect 1598 2808 1602 2812
rect 1646 2808 1650 2812
rect 1670 2808 1674 2812
rect 1774 2808 1778 2812
rect 2126 2808 2130 2812
rect 482 2803 486 2807
rect 490 2803 493 2807
rect 493 2803 494 2807
rect 1514 2803 1518 2807
rect 1522 2803 1525 2807
rect 1525 2803 1526 2807
rect 2538 2803 2542 2807
rect 2546 2803 2549 2807
rect 2549 2803 2550 2807
rect 470 2798 474 2802
rect 686 2798 690 2802
rect 814 2798 818 2802
rect 1806 2798 1810 2802
rect 1926 2798 1930 2802
rect 2182 2798 2186 2802
rect 2574 2798 2578 2802
rect 2590 2798 2594 2802
rect 566 2788 570 2792
rect 582 2788 586 2792
rect 806 2788 810 2792
rect 1110 2788 1114 2792
rect 1406 2788 1410 2792
rect 1542 2788 1546 2792
rect 2494 2788 2498 2792
rect 3454 2788 3458 2792
rect 262 2778 266 2782
rect 1046 2778 1050 2782
rect 1494 2778 1498 2782
rect 1726 2778 1730 2782
rect 1734 2778 1738 2782
rect 3478 2778 3482 2782
rect 950 2768 954 2772
rect 958 2768 962 2772
rect 1550 2768 1554 2772
rect 1790 2768 1794 2772
rect 1862 2768 1866 2772
rect 2102 2768 2106 2772
rect 2926 2768 2930 2772
rect 3022 2768 3026 2772
rect 3182 2768 3186 2772
rect 430 2758 434 2762
rect 854 2758 858 2762
rect 878 2758 882 2762
rect 1110 2758 1114 2762
rect 1254 2758 1258 2762
rect 1374 2758 1378 2762
rect 1454 2758 1458 2762
rect 1742 2758 1746 2762
rect 1950 2758 1954 2762
rect 2062 2758 2066 2762
rect 2166 2758 2170 2762
rect 2550 2758 2554 2762
rect 2734 2758 2738 2762
rect 3174 2758 3178 2762
rect 3198 2758 3202 2762
rect 334 2748 338 2752
rect 550 2748 554 2752
rect 870 2748 874 2752
rect 926 2748 930 2752
rect 950 2748 954 2752
rect 1086 2748 1090 2752
rect 1182 2748 1186 2752
rect 1198 2748 1202 2752
rect 1230 2748 1234 2752
rect 1238 2748 1242 2752
rect 1734 2748 1738 2752
rect 1846 2748 1850 2752
rect 2190 2748 2194 2752
rect 2286 2748 2290 2752
rect 2478 2748 2482 2752
rect 2638 2748 2642 2752
rect 2702 2748 2706 2752
rect 3230 2748 3234 2752
rect 3254 2748 3258 2752
rect 3542 2748 3546 2752
rect 38 2738 42 2742
rect 182 2738 186 2742
rect 534 2738 538 2742
rect 550 2738 554 2742
rect 878 2738 882 2742
rect 886 2738 890 2742
rect 1462 2738 1466 2742
rect 1966 2738 1970 2742
rect 478 2728 482 2732
rect 2070 2738 2074 2742
rect 2422 2738 2426 2742
rect 2486 2738 2490 2742
rect 2790 2738 2794 2742
rect 2838 2738 2842 2742
rect 2886 2738 2890 2742
rect 3382 2738 3386 2742
rect 3446 2738 3450 2742
rect 542 2728 546 2732
rect 646 2728 650 2732
rect 694 2728 698 2732
rect 1038 2728 1042 2732
rect 1110 2728 1114 2732
rect 1174 2728 1178 2732
rect 1366 2728 1370 2732
rect 1422 2728 1426 2732
rect 1574 2728 1578 2732
rect 1630 2728 1634 2732
rect 1726 2728 1730 2732
rect 2006 2728 2010 2732
rect 2086 2728 2090 2732
rect 2118 2728 2122 2732
rect 2134 2728 2138 2732
rect 2438 2728 2442 2732
rect 2798 2728 2802 2732
rect 3166 2728 3170 2732
rect 3318 2728 3322 2732
rect 286 2718 290 2722
rect 358 2718 362 2722
rect 1758 2718 1762 2722
rect 2118 2718 2122 2722
rect 2222 2718 2226 2722
rect 2526 2718 2530 2722
rect 2718 2718 2722 2722
rect 2934 2718 2938 2722
rect 2958 2718 2962 2722
rect 3030 2718 3034 2722
rect 3286 2718 3290 2722
rect 446 2708 450 2712
rect 494 2708 498 2712
rect 758 2708 762 2712
rect 1326 2708 1330 2712
rect 1358 2708 1362 2712
rect 1598 2708 1602 2712
rect 1790 2708 1794 2712
rect 2350 2708 2354 2712
rect 2590 2708 2594 2712
rect 994 2703 998 2707
rect 1002 2703 1005 2707
rect 1005 2703 1006 2707
rect 2026 2703 2030 2707
rect 2034 2703 2037 2707
rect 2037 2703 2038 2707
rect 3042 2703 3046 2707
rect 3050 2703 3053 2707
rect 3053 2703 3054 2707
rect 374 2698 378 2702
rect 454 2698 458 2702
rect 662 2698 666 2702
rect 718 2698 722 2702
rect 894 2698 898 2702
rect 918 2698 922 2702
rect 1038 2698 1042 2702
rect 1230 2698 1234 2702
rect 1918 2698 1922 2702
rect 1982 2698 1986 2702
rect 2342 2698 2346 2702
rect 2350 2698 2354 2702
rect 2654 2698 2658 2702
rect 2910 2698 2914 2702
rect 6 2688 10 2692
rect 406 2688 410 2692
rect 422 2688 426 2692
rect 446 2688 450 2692
rect 902 2688 906 2692
rect 1110 2688 1114 2692
rect 1670 2688 1674 2692
rect 1830 2688 1834 2692
rect 1998 2688 2002 2692
rect 2766 2688 2770 2692
rect 2814 2688 2818 2692
rect 3030 2688 3034 2692
rect 454 2678 458 2682
rect 566 2678 570 2682
rect 574 2678 578 2682
rect 742 2678 746 2682
rect 798 2678 802 2682
rect 1414 2678 1418 2682
rect 1734 2678 1738 2682
rect 2246 2678 2250 2682
rect 2310 2678 2314 2682
rect 2342 2678 2346 2682
rect 2366 2678 2370 2682
rect 2918 2678 2922 2682
rect 2990 2678 2994 2682
rect 3230 2678 3234 2682
rect 14 2668 18 2672
rect 22 2668 26 2672
rect 334 2668 338 2672
rect 1142 2668 1146 2672
rect 1158 2668 1162 2672
rect 1230 2668 1234 2672
rect 1470 2668 1474 2672
rect 1614 2668 1618 2672
rect 1902 2668 1906 2672
rect 1966 2668 1970 2672
rect 2126 2668 2130 2672
rect 2406 2668 2410 2672
rect 2414 2668 2418 2672
rect 230 2658 234 2662
rect 2590 2668 2594 2672
rect 2630 2668 2634 2672
rect 2734 2668 2738 2672
rect 2758 2668 2762 2672
rect 2822 2668 2826 2672
rect 3262 2668 3266 2672
rect 3334 2668 3338 2672
rect 510 2658 514 2662
rect 646 2658 650 2662
rect 950 2658 954 2662
rect 1054 2658 1058 2662
rect 1126 2658 1130 2662
rect 1446 2658 1450 2662
rect 1510 2658 1514 2662
rect 2118 2658 2122 2662
rect 2774 2658 2778 2662
rect 2830 2658 2834 2662
rect 2854 2658 2858 2662
rect 2990 2658 2994 2662
rect 3182 2658 3186 2662
rect 3270 2658 3274 2662
rect 6 2648 10 2652
rect 294 2648 298 2652
rect 334 2648 338 2652
rect 438 2648 442 2652
rect 558 2648 562 2652
rect 590 2648 594 2652
rect 774 2648 778 2652
rect 782 2648 786 2652
rect 1486 2648 1490 2652
rect 1638 2648 1642 2652
rect 1774 2648 1778 2652
rect 2054 2648 2058 2652
rect 2142 2648 2146 2652
rect 2638 2648 2642 2652
rect 3254 2648 3258 2652
rect 382 2638 386 2642
rect 542 2638 546 2642
rect 606 2638 610 2642
rect 646 2638 650 2642
rect 838 2638 842 2642
rect 950 2638 954 2642
rect 1646 2638 1650 2642
rect 1886 2638 1890 2642
rect 2158 2638 2162 2642
rect 2214 2638 2218 2642
rect 2646 2638 2650 2642
rect 2742 2638 2746 2642
rect 2766 2638 2770 2642
rect 2838 2638 2842 2642
rect 3318 2638 3322 2642
rect 22 2628 26 2632
rect 598 2628 602 2632
rect 862 2628 866 2632
rect 878 2628 882 2632
rect 910 2628 914 2632
rect 926 2628 930 2632
rect 974 2628 978 2632
rect 2790 2628 2794 2632
rect 2998 2628 3002 2632
rect 142 2618 146 2622
rect 350 2618 354 2622
rect 1678 2618 1682 2622
rect 1830 2618 1834 2622
rect 1910 2618 1914 2622
rect 1918 2618 1922 2622
rect 2494 2618 2498 2622
rect 2654 2618 2658 2622
rect 3222 2618 3226 2622
rect 3382 2618 3386 2622
rect 30 2608 34 2612
rect 574 2608 578 2612
rect 1054 2608 1058 2612
rect 1790 2608 1794 2612
rect 1878 2608 1882 2612
rect 2038 2608 2042 2612
rect 2510 2608 2514 2612
rect 2590 2608 2594 2612
rect 2934 2608 2938 2612
rect 482 2603 486 2607
rect 490 2603 493 2607
rect 493 2603 494 2607
rect 1514 2603 1518 2607
rect 1522 2603 1525 2607
rect 1525 2603 1526 2607
rect 2538 2603 2542 2607
rect 2546 2603 2549 2607
rect 2549 2603 2550 2607
rect 438 2598 442 2602
rect 846 2598 850 2602
rect 1174 2598 1178 2602
rect 1302 2598 1306 2602
rect 1478 2598 1482 2602
rect 1838 2598 1842 2602
rect 1862 2598 1866 2602
rect 2222 2598 2226 2602
rect 2558 2598 2562 2602
rect 3422 2598 3426 2602
rect 142 2588 146 2592
rect 454 2588 458 2592
rect 622 2588 626 2592
rect 1510 2588 1514 2592
rect 1798 2588 1802 2592
rect 1846 2588 1850 2592
rect 1870 2588 1874 2592
rect 3526 2588 3530 2592
rect 878 2578 882 2582
rect 894 2578 898 2582
rect 910 2578 914 2582
rect 1390 2578 1394 2582
rect 1758 2578 1762 2582
rect 2558 2578 2562 2582
rect 2606 2578 2610 2582
rect 2622 2578 2626 2582
rect 630 2568 634 2572
rect 1254 2568 1258 2572
rect 2006 2568 2010 2572
rect 2430 2568 2434 2572
rect 2974 2568 2978 2572
rect 326 2558 330 2562
rect 430 2558 434 2562
rect 614 2558 618 2562
rect 718 2558 722 2562
rect 766 2558 770 2562
rect 838 2558 842 2562
rect 1038 2558 1042 2562
rect 1086 2558 1090 2562
rect 1118 2558 1122 2562
rect 1454 2558 1458 2562
rect 1510 2558 1514 2562
rect 1694 2558 1698 2562
rect 1774 2558 1778 2562
rect 1822 2558 1826 2562
rect 2462 2558 2466 2562
rect 2526 2558 2530 2562
rect 2798 2558 2802 2562
rect 2950 2558 2954 2562
rect 6 2548 10 2552
rect 286 2548 290 2552
rect 534 2548 538 2552
rect 1174 2548 1178 2552
rect 1214 2548 1218 2552
rect 1430 2548 1434 2552
rect 1574 2548 1578 2552
rect 1670 2548 1674 2552
rect 1726 2548 1730 2552
rect 1734 2548 1738 2552
rect 2046 2548 2050 2552
rect 2318 2548 2322 2552
rect 2350 2548 2354 2552
rect 2774 2548 2778 2552
rect 2870 2548 2874 2552
rect 6 2538 10 2542
rect 582 2538 586 2542
rect 718 2538 722 2542
rect 918 2538 922 2542
rect 942 2538 946 2542
rect 1006 2538 1010 2542
rect 1030 2538 1034 2542
rect 1078 2538 1082 2542
rect 1142 2538 1146 2542
rect 1454 2538 1458 2542
rect 1782 2538 1786 2542
rect 1830 2538 1834 2542
rect 1894 2538 1898 2542
rect 1982 2538 1986 2542
rect 2070 2538 2074 2542
rect 30 2528 34 2532
rect 814 2528 818 2532
rect 998 2528 1002 2532
rect 1134 2528 1138 2532
rect 1278 2528 1282 2532
rect 1686 2528 1690 2532
rect 2406 2538 2410 2542
rect 2486 2538 2490 2542
rect 2590 2538 2594 2542
rect 2606 2538 2610 2542
rect 2846 2538 2850 2542
rect 3158 2538 3162 2542
rect 1918 2528 1922 2532
rect 2062 2528 2066 2532
rect 2182 2528 2186 2532
rect 2206 2528 2210 2532
rect 2254 2528 2258 2532
rect 2350 2528 2354 2532
rect 2470 2528 2474 2532
rect 2518 2528 2522 2532
rect 2534 2528 2538 2532
rect 3246 2528 3250 2532
rect 62 2518 66 2522
rect 150 2518 154 2522
rect 366 2518 370 2522
rect 430 2518 434 2522
rect 614 2518 618 2522
rect 774 2518 778 2522
rect 1062 2518 1066 2522
rect 1222 2518 1226 2522
rect 1358 2518 1362 2522
rect 1846 2518 1850 2522
rect 2382 2518 2386 2522
rect 2398 2518 2402 2522
rect 2430 2518 2434 2522
rect 2454 2518 2458 2522
rect 182 2508 186 2512
rect 814 2508 818 2512
rect 974 2508 978 2512
rect 1086 2508 1090 2512
rect 1118 2508 1122 2512
rect 1334 2508 1338 2512
rect 1406 2508 1410 2512
rect 1558 2508 1562 2512
rect 1622 2508 1626 2512
rect 1646 2508 1650 2512
rect 2414 2508 2418 2512
rect 3150 2508 3154 2512
rect 3166 2508 3170 2512
rect 994 2503 998 2507
rect 1002 2503 1005 2507
rect 1005 2503 1006 2507
rect 2026 2503 2030 2507
rect 2034 2503 2037 2507
rect 2037 2503 2038 2507
rect 3042 2503 3046 2507
rect 3050 2503 3053 2507
rect 3053 2503 3054 2507
rect 198 2498 202 2502
rect 214 2498 218 2502
rect 454 2498 458 2502
rect 462 2498 466 2502
rect 758 2498 762 2502
rect 806 2498 810 2502
rect 1014 2498 1018 2502
rect 1246 2498 1250 2502
rect 1334 2498 1338 2502
rect 1662 2498 1666 2502
rect 1734 2498 1738 2502
rect 2046 2498 2050 2502
rect 2134 2498 2138 2502
rect 86 2488 90 2492
rect 550 2488 554 2492
rect 598 2488 602 2492
rect 606 2488 610 2492
rect 1006 2488 1010 2492
rect 1062 2488 1066 2492
rect 1078 2488 1082 2492
rect 1254 2488 1258 2492
rect 1262 2488 1266 2492
rect 1374 2488 1378 2492
rect 1630 2488 1634 2492
rect 1654 2488 1658 2492
rect 1766 2488 1770 2492
rect 1790 2488 1794 2492
rect 1830 2488 1834 2492
rect 2006 2488 2010 2492
rect 2150 2488 2154 2492
rect 2326 2488 2330 2492
rect 2582 2488 2586 2492
rect 2598 2488 2602 2492
rect 2622 2488 2626 2492
rect 2726 2488 2730 2492
rect 2950 2488 2954 2492
rect 3126 2488 3130 2492
rect 318 2478 322 2482
rect 462 2478 466 2482
rect 686 2478 690 2482
rect 694 2478 698 2482
rect 1102 2478 1106 2482
rect 1406 2478 1410 2482
rect 1534 2478 1538 2482
rect 1678 2478 1682 2482
rect 2254 2478 2258 2482
rect 3334 2478 3338 2482
rect 3366 2478 3370 2482
rect 22 2468 26 2472
rect 302 2468 306 2472
rect 446 2468 450 2472
rect 806 2468 810 2472
rect 878 2468 882 2472
rect 926 2468 930 2472
rect 1038 2468 1042 2472
rect 1302 2468 1306 2472
rect 1382 2468 1386 2472
rect 1390 2468 1394 2472
rect 1486 2468 1490 2472
rect 1502 2468 1506 2472
rect 2006 2468 2010 2472
rect 2062 2468 2066 2472
rect 2366 2468 2370 2472
rect 2478 2468 2482 2472
rect 2830 2468 2834 2472
rect 3166 2468 3170 2472
rect 3174 2468 3178 2472
rect 3342 2468 3346 2472
rect 14 2458 18 2462
rect 574 2458 578 2462
rect 662 2458 666 2462
rect 670 2458 674 2462
rect 750 2458 754 2462
rect 838 2458 842 2462
rect 894 2458 898 2462
rect 1070 2458 1074 2462
rect 1246 2458 1250 2462
rect 1294 2458 1298 2462
rect 1398 2458 1402 2462
rect 2254 2458 2258 2462
rect 2294 2458 2298 2462
rect 2510 2458 2514 2462
rect 2550 2458 2554 2462
rect 2590 2458 2594 2462
rect 2782 2458 2786 2462
rect 2958 2458 2962 2462
rect 3254 2458 3258 2462
rect 3422 2458 3426 2462
rect 62 2448 66 2452
rect 694 2448 698 2452
rect 974 2448 978 2452
rect 1094 2448 1098 2452
rect 1110 2448 1114 2452
rect 1214 2448 1218 2452
rect 1286 2448 1290 2452
rect 1438 2448 1442 2452
rect 1526 2448 1530 2452
rect 1590 2448 1594 2452
rect 1734 2448 1738 2452
rect 2286 2448 2290 2452
rect 2470 2448 2474 2452
rect 2478 2448 2482 2452
rect 2958 2448 2962 2452
rect 3142 2448 3146 2452
rect 3190 2448 3194 2452
rect 3350 2448 3354 2452
rect 758 2438 762 2442
rect 870 2438 874 2442
rect 1014 2438 1018 2442
rect 1134 2438 1138 2442
rect 1190 2438 1194 2442
rect 1318 2438 1322 2442
rect 1398 2438 1402 2442
rect 2518 2438 2522 2442
rect 2774 2438 2778 2442
rect 3142 2438 3146 2442
rect 3534 2438 3538 2442
rect 158 2428 162 2432
rect 422 2428 426 2432
rect 510 2428 514 2432
rect 1182 2428 1186 2432
rect 2526 2428 2530 2432
rect 3158 2428 3162 2432
rect 3270 2428 3274 2432
rect 142 2418 146 2422
rect 694 2418 698 2422
rect 1574 2418 1578 2422
rect 1646 2418 1650 2422
rect 1982 2418 1986 2422
rect 2742 2418 2746 2422
rect 2886 2418 2890 2422
rect 2918 2418 2922 2422
rect 470 2408 474 2412
rect 846 2408 850 2412
rect 1198 2408 1202 2412
rect 1230 2408 1234 2412
rect 1366 2408 1370 2412
rect 1414 2408 1418 2412
rect 2198 2408 2202 2412
rect 2638 2408 2642 2412
rect 482 2403 486 2407
rect 490 2403 493 2407
rect 493 2403 494 2407
rect 6 2398 10 2402
rect 502 2398 506 2402
rect 686 2398 690 2402
rect 966 2398 970 2402
rect 1022 2398 1026 2402
rect 1054 2398 1058 2402
rect 1514 2403 1518 2407
rect 1522 2403 1525 2407
rect 1525 2403 1526 2407
rect 2538 2403 2542 2407
rect 2546 2403 2549 2407
rect 2549 2403 2550 2407
rect 1390 2398 1394 2402
rect 2046 2398 2050 2402
rect 2646 2398 2650 2402
rect 2854 2398 2858 2402
rect 3366 2398 3370 2402
rect 438 2388 442 2392
rect 878 2388 882 2392
rect 1646 2388 1650 2392
rect 2398 2388 2402 2392
rect 3134 2388 3138 2392
rect 518 2378 522 2382
rect 638 2378 642 2382
rect 766 2378 770 2382
rect 1142 2378 1146 2382
rect 1166 2378 1170 2382
rect 2854 2378 2858 2382
rect 6 2368 10 2372
rect 294 2368 298 2372
rect 334 2368 338 2372
rect 350 2368 354 2372
rect 582 2368 586 2372
rect 758 2368 762 2372
rect 814 2368 818 2372
rect 1070 2368 1074 2372
rect 1134 2368 1138 2372
rect 1294 2368 1298 2372
rect 1446 2368 1450 2372
rect 1878 2368 1882 2372
rect 1894 2368 1898 2372
rect 2366 2368 2370 2372
rect 2686 2368 2690 2372
rect 2766 2368 2770 2372
rect 718 2358 722 2362
rect 830 2358 834 2362
rect 878 2358 882 2362
rect 1022 2358 1026 2362
rect 1038 2358 1042 2362
rect 1582 2358 1586 2362
rect 2126 2358 2130 2362
rect 2470 2358 2474 2362
rect 2582 2358 2586 2362
rect 2590 2358 2594 2362
rect 2942 2358 2946 2362
rect 2950 2358 2954 2362
rect 2974 2358 2978 2362
rect 3198 2358 3202 2362
rect 3350 2358 3354 2362
rect 3406 2358 3410 2362
rect 6 2348 10 2352
rect 542 2348 546 2352
rect 622 2348 626 2352
rect 654 2348 658 2352
rect 702 2348 706 2352
rect 710 2348 714 2352
rect 790 2348 794 2352
rect 886 2348 890 2352
rect 918 2348 922 2352
rect 934 2348 938 2352
rect 1046 2348 1050 2352
rect 1062 2348 1066 2352
rect 1246 2348 1250 2352
rect 1270 2348 1274 2352
rect 1358 2348 1362 2352
rect 1414 2348 1418 2352
rect 1646 2348 1650 2352
rect 1662 2348 1666 2352
rect 1998 2348 2002 2352
rect 2094 2348 2098 2352
rect 2110 2348 2114 2352
rect 2230 2348 2234 2352
rect 2334 2348 2338 2352
rect 2422 2348 2426 2352
rect 2486 2348 2490 2352
rect 2702 2348 2706 2352
rect 3206 2348 3210 2352
rect 3334 2348 3338 2352
rect 30 2338 34 2342
rect 390 2338 394 2342
rect 414 2338 418 2342
rect 542 2338 546 2342
rect 558 2338 562 2342
rect 662 2338 666 2342
rect 782 2338 786 2342
rect 814 2338 818 2342
rect 918 2338 922 2342
rect 1142 2338 1146 2342
rect 1166 2338 1170 2342
rect 1214 2338 1218 2342
rect 1254 2338 1258 2342
rect 1334 2338 1338 2342
rect 1406 2338 1410 2342
rect 1502 2338 1506 2342
rect 1726 2338 1730 2342
rect 1742 2338 1746 2342
rect 1774 2338 1778 2342
rect 1942 2338 1946 2342
rect 2270 2338 2274 2342
rect 2774 2338 2778 2342
rect 2862 2338 2866 2342
rect 2926 2338 2930 2342
rect 3118 2338 3122 2342
rect 3366 2338 3370 2342
rect 3382 2338 3386 2342
rect 3446 2338 3450 2342
rect 3462 2338 3466 2342
rect 174 2328 178 2332
rect 182 2328 186 2332
rect 342 2328 346 2332
rect 374 2328 378 2332
rect 534 2328 538 2332
rect 870 2328 874 2332
rect 1134 2328 1138 2332
rect 1518 2328 1522 2332
rect 1710 2328 1714 2332
rect 1742 2328 1746 2332
rect 1782 2328 1786 2332
rect 1838 2328 1842 2332
rect 1950 2328 1954 2332
rect 2006 2328 2010 2332
rect 2094 2328 2098 2332
rect 2446 2328 2450 2332
rect 2510 2328 2514 2332
rect 2558 2328 2562 2332
rect 2582 2328 2586 2332
rect 2950 2328 2954 2332
rect 3318 2328 3322 2332
rect 550 2318 554 2322
rect 574 2318 578 2322
rect 598 2318 602 2322
rect 718 2318 722 2322
rect 742 2318 746 2322
rect 782 2318 786 2322
rect 862 2318 866 2322
rect 2014 2318 2018 2322
rect 2678 2318 2682 2322
rect 2694 2318 2698 2322
rect 2966 2318 2970 2322
rect 2974 2318 2978 2322
rect 3278 2318 3282 2322
rect 422 2308 426 2312
rect 966 2308 970 2312
rect 1150 2308 1154 2312
rect 1206 2308 1210 2312
rect 1214 2308 1218 2312
rect 1286 2308 1290 2312
rect 1838 2308 1842 2312
rect 2758 2308 2762 2312
rect 2902 2308 2906 2312
rect 3382 2308 3386 2312
rect 994 2303 998 2307
rect 1002 2303 1005 2307
rect 1005 2303 1006 2307
rect 558 2298 562 2302
rect 982 2298 986 2302
rect 1014 2298 1018 2302
rect 1278 2298 1282 2302
rect 1758 2298 1762 2302
rect 2026 2303 2030 2307
rect 2034 2303 2037 2307
rect 2037 2303 2038 2307
rect 2638 2298 2642 2302
rect 2670 2298 2674 2302
rect 3042 2303 3046 2307
rect 3050 2303 3053 2307
rect 3053 2303 3054 2307
rect 2918 2298 2922 2302
rect 454 2288 458 2292
rect 1118 2288 1122 2292
rect 1150 2288 1154 2292
rect 1238 2288 1242 2292
rect 1262 2288 1266 2292
rect 1430 2288 1434 2292
rect 1542 2288 1546 2292
rect 1894 2288 1898 2292
rect 1958 2288 1962 2292
rect 2326 2288 2330 2292
rect 2438 2288 2442 2292
rect 3102 2288 3106 2292
rect 3134 2288 3138 2292
rect 3206 2288 3210 2292
rect 3326 2288 3330 2292
rect 3366 2288 3370 2292
rect 3422 2288 3426 2292
rect 606 2278 610 2282
rect 718 2278 722 2282
rect 902 2278 906 2282
rect 958 2278 962 2282
rect 1038 2278 1042 2282
rect 1062 2278 1066 2282
rect 1118 2278 1122 2282
rect 1134 2278 1138 2282
rect 1190 2278 1194 2282
rect 1222 2278 1226 2282
rect 1278 2278 1282 2282
rect 1294 2278 1298 2282
rect 1430 2278 1434 2282
rect 1454 2278 1458 2282
rect 1686 2278 1690 2282
rect 1726 2278 1730 2282
rect 1966 2278 1970 2282
rect 2110 2278 2114 2282
rect 2150 2278 2154 2282
rect 2430 2278 2434 2282
rect 2462 2278 2466 2282
rect 2582 2278 2586 2282
rect 2598 2278 2602 2282
rect 3150 2278 3154 2282
rect 6 2268 10 2272
rect 78 2268 82 2272
rect 102 2268 106 2272
rect 342 2268 346 2272
rect 358 2268 362 2272
rect 430 2268 434 2272
rect 758 2268 762 2272
rect 846 2268 850 2272
rect 886 2268 890 2272
rect 894 2268 898 2272
rect 1246 2268 1250 2272
rect 1310 2268 1314 2272
rect 1534 2268 1538 2272
rect 1574 2268 1578 2272
rect 1622 2268 1626 2272
rect 1694 2268 1698 2272
rect 2014 2268 2018 2272
rect 2070 2268 2074 2272
rect 2126 2268 2130 2272
rect 2134 2268 2138 2272
rect 2166 2268 2170 2272
rect 2190 2268 2194 2272
rect 2206 2268 2210 2272
rect 2478 2268 2482 2272
rect 2486 2268 2490 2272
rect 3206 2268 3210 2272
rect 806 2258 810 2262
rect 1094 2258 1098 2262
rect 1142 2258 1146 2262
rect 1910 2258 1914 2262
rect 2022 2258 2026 2262
rect 14 2248 18 2252
rect 566 2248 570 2252
rect 582 2248 586 2252
rect 734 2248 738 2252
rect 742 2248 746 2252
rect 1158 2248 1162 2252
rect 1166 2248 1170 2252
rect 1702 2248 1706 2252
rect 1710 2248 1714 2252
rect 2302 2248 2306 2252
rect 2406 2248 2410 2252
rect 2518 2248 2522 2252
rect 2638 2248 2642 2252
rect 2854 2248 2858 2252
rect 2870 2248 2874 2252
rect 3086 2248 3090 2252
rect 3238 2248 3242 2252
rect 38 2238 42 2242
rect 510 2238 514 2242
rect 526 2238 530 2242
rect 638 2238 642 2242
rect 678 2238 682 2242
rect 758 2238 762 2242
rect 870 2238 874 2242
rect 1638 2238 1642 2242
rect 2502 2238 2506 2242
rect 2566 2238 2570 2242
rect 3246 2238 3250 2242
rect 6 2228 10 2232
rect 1174 2228 1178 2232
rect 1582 2228 1586 2232
rect 2174 2228 2178 2232
rect 3294 2228 3298 2232
rect 502 2218 506 2222
rect 1110 2218 1114 2222
rect 1126 2218 1130 2222
rect 1654 2218 1658 2222
rect 2806 2218 2810 2222
rect 2990 2218 2994 2222
rect 2998 2218 3002 2222
rect 3190 2218 3194 2222
rect 3238 2218 3242 2222
rect 3342 2218 3346 2222
rect 286 2208 290 2212
rect 590 2208 594 2212
rect 2510 2208 2514 2212
rect 2766 2208 2770 2212
rect 482 2203 486 2207
rect 490 2203 493 2207
rect 493 2203 494 2207
rect 1514 2203 1518 2207
rect 1522 2203 1525 2207
rect 1525 2203 1526 2207
rect 2538 2203 2542 2207
rect 2546 2203 2549 2207
rect 2549 2203 2550 2207
rect 238 2198 242 2202
rect 366 2198 370 2202
rect 502 2198 506 2202
rect 814 2198 818 2202
rect 1086 2198 1090 2202
rect 1454 2198 1458 2202
rect 1542 2198 1546 2202
rect 1790 2198 1794 2202
rect 1806 2198 1810 2202
rect 1886 2198 1890 2202
rect 2062 2198 2066 2202
rect 2070 2198 2074 2202
rect 2086 2198 2090 2202
rect 2798 2198 2802 2202
rect 958 2188 962 2192
rect 1374 2188 1378 2192
rect 134 2178 138 2182
rect 1422 2178 1426 2182
rect 1542 2178 1546 2182
rect 1550 2178 1554 2182
rect 1718 2178 1722 2182
rect 1902 2178 1906 2182
rect 1910 2178 1914 2182
rect 22 2168 26 2172
rect 318 2168 322 2172
rect 374 2168 378 2172
rect 630 2168 634 2172
rect 686 2168 690 2172
rect 702 2168 706 2172
rect 822 2168 826 2172
rect 862 2168 866 2172
rect 902 2168 906 2172
rect 950 2168 954 2172
rect 990 2168 994 2172
rect 2054 2168 2058 2172
rect 2086 2168 2090 2172
rect 2102 2168 2106 2172
rect 2238 2168 2242 2172
rect 2382 2168 2386 2172
rect 2686 2168 2690 2172
rect 3454 2168 3458 2172
rect 278 2158 282 2162
rect 502 2158 506 2162
rect 542 2158 546 2162
rect 558 2158 562 2162
rect 582 2158 586 2162
rect 790 2158 794 2162
rect 2094 2158 2098 2162
rect 2254 2158 2258 2162
rect 2366 2158 2370 2162
rect 2470 2158 2474 2162
rect 2910 2158 2914 2162
rect 2934 2158 2938 2162
rect 166 2148 170 2152
rect 230 2148 234 2152
rect 606 2148 610 2152
rect 902 2148 906 2152
rect 1014 2148 1018 2152
rect 1142 2148 1146 2152
rect 1294 2148 1298 2152
rect 1630 2148 1634 2152
rect 2094 2148 2098 2152
rect 3158 2148 3162 2152
rect 3198 2148 3202 2152
rect 3222 2148 3226 2152
rect 3342 2148 3346 2152
rect 3446 2148 3450 2152
rect 174 2138 178 2142
rect 558 2138 562 2142
rect 574 2138 578 2142
rect 774 2138 778 2142
rect 798 2138 802 2142
rect 998 2138 1002 2142
rect 1126 2138 1130 2142
rect 1158 2138 1162 2142
rect 1646 2138 1650 2142
rect 1790 2138 1794 2142
rect 1822 2138 1826 2142
rect 1838 2138 1842 2142
rect 1958 2138 1962 2142
rect 2494 2138 2498 2142
rect 2534 2138 2538 2142
rect 2646 2138 2650 2142
rect 3486 2138 3490 2142
rect 190 2128 194 2132
rect 310 2128 314 2132
rect 342 2128 346 2132
rect 646 2128 650 2132
rect 982 2128 986 2132
rect 1294 2128 1298 2132
rect 1790 2128 1794 2132
rect 1814 2128 1818 2132
rect 1918 2128 1922 2132
rect 2238 2128 2242 2132
rect 2574 2128 2578 2132
rect 3294 2128 3298 2132
rect 3342 2128 3346 2132
rect 550 2118 554 2122
rect 1102 2118 1106 2122
rect 1206 2118 1210 2122
rect 1254 2118 1258 2122
rect 1894 2118 1898 2122
rect 2830 2118 2834 2122
rect 630 2108 634 2112
rect 1286 2108 1290 2112
rect 1862 2108 1866 2112
rect 2046 2108 2050 2112
rect 2182 2108 2186 2112
rect 2286 2108 2290 2112
rect 2358 2108 2362 2112
rect 2742 2108 2746 2112
rect 2910 2108 2914 2112
rect 3238 2108 3242 2112
rect 3262 2108 3266 2112
rect 3446 2108 3450 2112
rect 994 2103 998 2107
rect 1002 2103 1005 2107
rect 1005 2103 1006 2107
rect 238 2098 242 2102
rect 750 2098 754 2102
rect 1334 2098 1338 2102
rect 1462 2098 1466 2102
rect 2026 2103 2030 2107
rect 2034 2103 2037 2107
rect 2037 2103 2038 2107
rect 3042 2103 3046 2107
rect 3050 2103 3053 2107
rect 3053 2103 3054 2107
rect 1646 2098 1650 2102
rect 1750 2098 1754 2102
rect 1846 2098 1850 2102
rect 1854 2098 1858 2102
rect 2214 2098 2218 2102
rect 2342 2098 2346 2102
rect 2478 2098 2482 2102
rect 3030 2098 3034 2102
rect 3486 2098 3490 2102
rect 182 2088 186 2092
rect 526 2088 530 2092
rect 782 2088 786 2092
rect 822 2088 826 2092
rect 910 2088 914 2092
rect 1046 2088 1050 2092
rect 1198 2088 1202 2092
rect 262 2078 266 2082
rect 318 2078 322 2082
rect 630 2078 634 2082
rect 694 2078 698 2082
rect 934 2078 938 2082
rect 1062 2078 1066 2082
rect 1262 2078 1266 2082
rect 1390 2078 1394 2082
rect 1494 2078 1498 2082
rect 1614 2078 1618 2082
rect 1766 2078 1770 2082
rect 1822 2078 1826 2082
rect 1910 2078 1914 2082
rect 2062 2078 2066 2082
rect 2150 2078 2154 2082
rect 2166 2078 2170 2082
rect 2206 2078 2210 2082
rect 2222 2078 2226 2082
rect 2342 2078 2346 2082
rect 2398 2078 2402 2082
rect 2414 2078 2418 2082
rect 2446 2078 2450 2082
rect 2942 2078 2946 2082
rect 3134 2078 3138 2082
rect 86 2068 90 2072
rect 270 2068 274 2072
rect 534 2068 538 2072
rect 550 2068 554 2072
rect 622 2068 626 2072
rect 798 2068 802 2072
rect 926 2068 930 2072
rect 1310 2068 1314 2072
rect 1710 2068 1714 2072
rect 1726 2068 1730 2072
rect 1774 2068 1778 2072
rect 1886 2068 1890 2072
rect 1926 2068 1930 2072
rect 2294 2068 2298 2072
rect 2382 2068 2386 2072
rect 2742 2068 2746 2072
rect 2774 2068 2778 2072
rect 3150 2068 3154 2072
rect 3198 2068 3202 2072
rect 3238 2068 3242 2072
rect 3558 2068 3562 2072
rect 70 2058 74 2062
rect 142 2058 146 2062
rect 1062 2058 1066 2062
rect 1094 2058 1098 2062
rect 1694 2058 1698 2062
rect 1766 2058 1770 2062
rect 1878 2058 1882 2062
rect 2086 2058 2090 2062
rect 2094 2058 2098 2062
rect 2142 2058 2146 2062
rect 2190 2058 2194 2062
rect 2302 2058 2306 2062
rect 2318 2058 2322 2062
rect 2390 2058 2394 2062
rect 2486 2058 2490 2062
rect 2782 2058 2786 2062
rect 22 2048 26 2052
rect 758 2048 762 2052
rect 910 2048 914 2052
rect 950 2048 954 2052
rect 1502 2048 1506 2052
rect 1574 2048 1578 2052
rect 1630 2048 1634 2052
rect 1854 2048 1858 2052
rect 1894 2048 1898 2052
rect 1998 2048 2002 2052
rect 2062 2048 2066 2052
rect 2134 2048 2138 2052
rect 2262 2048 2266 2052
rect 2342 2048 2346 2052
rect 2398 2048 2402 2052
rect 2414 2048 2418 2052
rect 2654 2048 2658 2052
rect 2718 2048 2722 2052
rect 2902 2048 2906 2052
rect 3038 2048 3042 2052
rect 3358 2048 3362 2052
rect 606 2038 610 2042
rect 710 2038 714 2042
rect 830 2038 834 2042
rect 1030 2038 1034 2042
rect 1254 2038 1258 2042
rect 1278 2038 1282 2042
rect 2198 2038 2202 2042
rect 2310 2038 2314 2042
rect 2486 2038 2490 2042
rect 2590 2038 2594 2042
rect 2790 2038 2794 2042
rect 3014 2038 3018 2042
rect 3126 2038 3130 2042
rect 302 2028 306 2032
rect 510 2028 514 2032
rect 838 2028 842 2032
rect 1022 2028 1026 2032
rect 1086 2028 1090 2032
rect 1414 2028 1418 2032
rect 1606 2028 1610 2032
rect 1734 2028 1738 2032
rect 1750 2028 1754 2032
rect 1838 2028 1842 2032
rect 2878 2028 2882 2032
rect 1662 2018 1666 2022
rect 1774 2018 1778 2022
rect 1934 2018 1938 2022
rect 1942 2018 1946 2022
rect 1958 2018 1962 2022
rect 2654 2018 2658 2022
rect 2918 2018 2922 2022
rect 174 2008 178 2012
rect 430 2008 434 2012
rect 942 2008 946 2012
rect 1598 2008 1602 2012
rect 1702 2008 1706 2012
rect 1918 2008 1922 2012
rect 1950 2008 1954 2012
rect 2438 2008 2442 2012
rect 2510 2008 2514 2012
rect 2886 2008 2890 2012
rect 3118 2008 3122 2012
rect 482 2003 486 2007
rect 490 2003 493 2007
rect 493 2003 494 2007
rect 1514 2003 1518 2007
rect 1522 2003 1525 2007
rect 1525 2003 1526 2007
rect 2538 2003 2542 2007
rect 2546 2003 2549 2007
rect 2549 2003 2550 2007
rect 462 1998 466 2002
rect 542 1998 546 2002
rect 1310 1998 1314 2002
rect 1342 1998 1346 2002
rect 1438 1998 1442 2002
rect 1542 1998 1546 2002
rect 1606 1998 1610 2002
rect 1662 1998 1666 2002
rect 1710 1998 1714 2002
rect 1926 1998 1930 2002
rect 1934 1998 1938 2002
rect 2142 1998 2146 2002
rect 2430 1998 2434 2002
rect 2446 1998 2450 2002
rect 2678 1998 2682 2002
rect 2894 1998 2898 2002
rect 358 1988 362 1992
rect 470 1988 474 1992
rect 582 1988 586 1992
rect 646 1988 650 1992
rect 654 1988 658 1992
rect 670 1988 674 1992
rect 774 1988 778 1992
rect 798 1988 802 1992
rect 886 1988 890 1992
rect 958 1988 962 1992
rect 1166 1988 1170 1992
rect 1294 1988 1298 1992
rect 2734 1988 2738 1992
rect 2750 1988 2754 1992
rect 2870 1988 2874 1992
rect 2926 1988 2930 1992
rect 3414 1988 3418 1992
rect 166 1978 170 1982
rect 318 1978 322 1982
rect 414 1978 418 1982
rect 438 1978 442 1982
rect 526 1978 530 1982
rect 726 1978 730 1982
rect 766 1978 770 1982
rect 1150 1978 1154 1982
rect 1774 1978 1778 1982
rect 1830 1978 1834 1982
rect 1998 1978 2002 1982
rect 2694 1978 2698 1982
rect 2878 1978 2882 1982
rect 566 1968 570 1972
rect 1046 1968 1050 1972
rect 1118 1968 1122 1972
rect 1246 1968 1250 1972
rect 1478 1968 1482 1972
rect 1726 1968 1730 1972
rect 1862 1968 1866 1972
rect 2046 1968 2050 1972
rect 2094 1968 2098 1972
rect 2206 1968 2210 1972
rect 2278 1968 2282 1972
rect 3006 1968 3010 1972
rect 118 1958 122 1962
rect 158 1958 162 1962
rect 462 1958 466 1962
rect 606 1958 610 1962
rect 638 1958 642 1962
rect 678 1958 682 1962
rect 1342 1958 1346 1962
rect 1358 1958 1362 1962
rect 1462 1958 1466 1962
rect 1486 1958 1490 1962
rect 1590 1958 1594 1962
rect 1662 1958 1666 1962
rect 1718 1958 1722 1962
rect 1822 1958 1826 1962
rect 1926 1958 1930 1962
rect 2270 1958 2274 1962
rect 2686 1958 2690 1962
rect 2926 1958 2930 1962
rect 3198 1958 3202 1962
rect 3262 1958 3266 1962
rect 3278 1958 3282 1962
rect 3334 1958 3338 1962
rect 3342 1958 3346 1962
rect 134 1948 138 1952
rect 214 1948 218 1952
rect 286 1948 290 1952
rect 430 1948 434 1952
rect 614 1948 618 1952
rect 902 1948 906 1952
rect 1134 1948 1138 1952
rect 1182 1948 1186 1952
rect 1302 1948 1306 1952
rect 1326 1948 1330 1952
rect 1406 1948 1410 1952
rect 1438 1948 1442 1952
rect 1670 1948 1674 1952
rect 1774 1948 1778 1952
rect 1782 1948 1786 1952
rect 1854 1948 1858 1952
rect 2006 1948 2010 1952
rect 2382 1948 2386 1952
rect 2478 1948 2482 1952
rect 2606 1948 2610 1952
rect 2766 1948 2770 1952
rect 2918 1948 2922 1952
rect 3270 1948 3274 1952
rect 526 1938 530 1942
rect 942 1938 946 1942
rect 982 1938 986 1942
rect 1254 1938 1258 1942
rect 1286 1938 1290 1942
rect 1430 1938 1434 1942
rect 1550 1938 1554 1942
rect 1574 1938 1578 1942
rect 1622 1938 1626 1942
rect 1742 1938 1746 1942
rect 1758 1938 1762 1942
rect 2094 1938 2098 1942
rect 2310 1938 2314 1942
rect 2526 1938 2530 1942
rect 2702 1938 2706 1942
rect 2910 1938 2914 1942
rect 2934 1938 2938 1942
rect 2958 1938 2962 1942
rect 3054 1938 3058 1942
rect 3198 1938 3202 1942
rect 542 1928 546 1932
rect 678 1928 682 1932
rect 766 1928 770 1932
rect 1302 1928 1306 1932
rect 1390 1928 1394 1932
rect 1534 1928 1538 1932
rect 1566 1928 1570 1932
rect 1630 1928 1634 1932
rect 1742 1928 1746 1932
rect 1774 1928 1778 1932
rect 1806 1928 1810 1932
rect 1870 1928 1874 1932
rect 1886 1928 1890 1932
rect 1918 1928 1922 1932
rect 1942 1928 1946 1932
rect 1974 1928 1978 1932
rect 2374 1928 2378 1932
rect 2478 1928 2482 1932
rect 2950 1928 2954 1932
rect 3222 1928 3226 1932
rect 3270 1928 3274 1932
rect 102 1918 106 1922
rect 286 1918 290 1922
rect 1766 1918 1770 1922
rect 1838 1918 1842 1922
rect 1846 1918 1850 1922
rect 1862 1918 1866 1922
rect 2038 1918 2042 1922
rect 2238 1918 2242 1922
rect 2734 1918 2738 1922
rect 3278 1918 3282 1922
rect 222 1908 226 1912
rect 310 1908 314 1912
rect 694 1908 698 1912
rect 1054 1908 1058 1912
rect 1798 1908 1802 1912
rect 1990 1908 1994 1912
rect 2046 1908 2050 1912
rect 2150 1908 2154 1912
rect 2166 1908 2170 1912
rect 2486 1908 2490 1912
rect 2710 1908 2714 1912
rect 2758 1908 2762 1912
rect 2918 1908 2922 1912
rect 3214 1908 3218 1912
rect 994 1903 998 1907
rect 1002 1903 1005 1907
rect 1005 1903 1006 1907
rect 2026 1903 2030 1907
rect 2034 1903 2037 1907
rect 2037 1903 2038 1907
rect 3042 1903 3046 1907
rect 3050 1903 3053 1907
rect 3053 1903 3054 1907
rect 198 1898 202 1902
rect 422 1898 426 1902
rect 638 1898 642 1902
rect 686 1898 690 1902
rect 742 1898 746 1902
rect 926 1898 930 1902
rect 2158 1898 2162 1902
rect 2222 1898 2226 1902
rect 2622 1898 2626 1902
rect 2974 1898 2978 1902
rect 3502 1898 3506 1902
rect 3526 1898 3530 1902
rect 1286 1888 1290 1892
rect 2214 1888 2218 1892
rect 2230 1888 2234 1892
rect 2254 1888 2258 1892
rect 2302 1888 2306 1892
rect 2318 1888 2322 1892
rect 2486 1888 2490 1892
rect 3078 1888 3082 1892
rect 3126 1888 3130 1892
rect 3230 1888 3234 1892
rect 222 1878 226 1882
rect 510 1878 514 1882
rect 630 1878 634 1882
rect 638 1878 642 1882
rect 998 1878 1002 1882
rect 1094 1878 1098 1882
rect 1158 1878 1162 1882
rect 1502 1878 1506 1882
rect 1654 1878 1658 1882
rect 1926 1878 1930 1882
rect 2678 1878 2682 1882
rect 2686 1878 2690 1882
rect 2838 1878 2842 1882
rect 2918 1878 2922 1882
rect 110 1868 114 1872
rect 614 1868 618 1872
rect 998 1868 1002 1872
rect 1214 1868 1218 1872
rect 1278 1868 1282 1872
rect 1318 1868 1322 1872
rect 1374 1868 1378 1872
rect 1438 1868 1442 1872
rect 1454 1868 1458 1872
rect 1590 1868 1594 1872
rect 1662 1868 1666 1872
rect 1670 1868 1674 1872
rect 1886 1868 1890 1872
rect 2342 1868 2346 1872
rect 2382 1868 2386 1872
rect 2630 1868 2634 1872
rect 2710 1868 2714 1872
rect 2966 1868 2970 1872
rect 3006 1868 3010 1872
rect 3078 1868 3082 1872
rect 3254 1868 3258 1872
rect 3542 1868 3546 1872
rect 30 1858 34 1862
rect 230 1858 234 1862
rect 334 1858 338 1862
rect 582 1858 586 1862
rect 622 1858 626 1862
rect 926 1858 930 1862
rect 1398 1858 1402 1862
rect 1446 1858 1450 1862
rect 1494 1858 1498 1862
rect 1622 1858 1626 1862
rect 1638 1858 1642 1862
rect 1686 1858 1690 1862
rect 1702 1858 1706 1862
rect 1734 1858 1738 1862
rect 1758 1858 1762 1862
rect 1926 1858 1930 1862
rect 2158 1858 2162 1862
rect 2270 1858 2274 1862
rect 2286 1858 2290 1862
rect 2838 1858 2842 1862
rect 2998 1858 3002 1862
rect 3014 1858 3018 1862
rect 3126 1858 3130 1862
rect 102 1848 106 1852
rect 166 1848 170 1852
rect 446 1848 450 1852
rect 518 1848 522 1852
rect 526 1848 530 1852
rect 774 1848 778 1852
rect 958 1848 962 1852
rect 1342 1848 1346 1852
rect 1350 1848 1354 1852
rect 1454 1848 1458 1852
rect 1542 1848 1546 1852
rect 1598 1848 1602 1852
rect 1718 1848 1722 1852
rect 1806 1848 1810 1852
rect 1830 1848 1834 1852
rect 1870 1848 1874 1852
rect 1886 1848 1890 1852
rect 1894 1848 1898 1852
rect 1910 1848 1914 1852
rect 1990 1848 1994 1852
rect 2006 1848 2010 1852
rect 2022 1848 2026 1852
rect 2078 1848 2082 1852
rect 2286 1848 2290 1852
rect 2334 1848 2338 1852
rect 2582 1848 2586 1852
rect 3118 1848 3122 1852
rect 3150 1848 3154 1852
rect 590 1838 594 1842
rect 1142 1838 1146 1842
rect 1222 1838 1226 1842
rect 1398 1838 1402 1842
rect 1598 1838 1602 1842
rect 1606 1838 1610 1842
rect 2070 1838 2074 1842
rect 3542 1838 3546 1842
rect 126 1828 130 1832
rect 310 1828 314 1832
rect 358 1828 362 1832
rect 926 1828 930 1832
rect 1214 1828 1218 1832
rect 1630 1828 1634 1832
rect 1894 1828 1898 1832
rect 1918 1828 1922 1832
rect 1934 1828 1938 1832
rect 2270 1828 2274 1832
rect 2334 1828 2338 1832
rect 2614 1828 2618 1832
rect 2646 1828 2650 1832
rect 438 1818 442 1822
rect 974 1818 978 1822
rect 1294 1818 1298 1822
rect 1526 1818 1530 1822
rect 1606 1818 1610 1822
rect 2438 1818 2442 1822
rect 2558 1818 2562 1822
rect 2718 1818 2722 1822
rect 2934 1818 2938 1822
rect 3142 1818 3146 1822
rect 3326 1818 3330 1822
rect 326 1808 330 1812
rect 646 1808 650 1812
rect 1094 1808 1098 1812
rect 1278 1808 1282 1812
rect 1414 1808 1418 1812
rect 1422 1808 1426 1812
rect 1470 1808 1474 1812
rect 1542 1808 1546 1812
rect 1766 1808 1770 1812
rect 1782 1808 1786 1812
rect 1870 1808 1874 1812
rect 1926 1808 1930 1812
rect 1934 1808 1938 1812
rect 2422 1808 2426 1812
rect 2678 1808 2682 1812
rect 482 1803 486 1807
rect 490 1803 493 1807
rect 493 1803 494 1807
rect 1514 1803 1518 1807
rect 1522 1803 1525 1807
rect 1525 1803 1526 1807
rect 294 1798 298 1802
rect 406 1798 410 1802
rect 502 1798 506 1802
rect 830 1798 834 1802
rect 1078 1798 1082 1802
rect 1134 1798 1138 1802
rect 1182 1798 1186 1802
rect 1270 1798 1274 1802
rect 1326 1798 1330 1802
rect 1334 1798 1338 1802
rect 1470 1798 1474 1802
rect 1574 1798 1578 1802
rect 1670 1798 1674 1802
rect 1990 1798 1994 1802
rect 2070 1798 2074 1802
rect 2538 1803 2542 1807
rect 2546 1803 2549 1807
rect 2549 1803 2550 1807
rect 2494 1798 2498 1802
rect 2582 1798 2586 1802
rect 2766 1798 2770 1802
rect 958 1788 962 1792
rect 2198 1788 2202 1792
rect 2262 1788 2266 1792
rect 2278 1788 2282 1792
rect 2606 1788 2610 1792
rect 2654 1788 2658 1792
rect 2678 1788 2682 1792
rect 2934 1788 2938 1792
rect 3302 1788 3306 1792
rect 3390 1788 3394 1792
rect 254 1778 258 1782
rect 526 1778 530 1782
rect 910 1778 914 1782
rect 1062 1778 1066 1782
rect 1126 1778 1130 1782
rect 1254 1778 1258 1782
rect 1494 1778 1498 1782
rect 1502 1778 1506 1782
rect 1558 1778 1562 1782
rect 1718 1778 1722 1782
rect 1742 1778 1746 1782
rect 1926 1778 1930 1782
rect 1958 1778 1962 1782
rect 2790 1778 2794 1782
rect 3430 1778 3434 1782
rect 3558 1778 3562 1782
rect 166 1768 170 1772
rect 206 1768 210 1772
rect 262 1768 266 1772
rect 414 1768 418 1772
rect 686 1768 690 1772
rect 702 1768 706 1772
rect 774 1768 778 1772
rect 982 1768 986 1772
rect 1134 1768 1138 1772
rect 1326 1768 1330 1772
rect 1334 1768 1338 1772
rect 1710 1768 1714 1772
rect 1830 1768 1834 1772
rect 1870 1768 1874 1772
rect 1878 1768 1882 1772
rect 1918 1768 1922 1772
rect 2654 1768 2658 1772
rect 2830 1768 2834 1772
rect 3422 1768 3426 1772
rect 134 1758 138 1762
rect 710 1758 714 1762
rect 726 1758 730 1762
rect 1046 1758 1050 1762
rect 1150 1758 1154 1762
rect 1254 1758 1258 1762
rect 1350 1758 1354 1762
rect 1438 1758 1442 1762
rect 1494 1758 1498 1762
rect 1582 1758 1586 1762
rect 1750 1758 1754 1762
rect 1854 1758 1858 1762
rect 1942 1758 1946 1762
rect 1958 1758 1962 1762
rect 2110 1758 2114 1762
rect 2286 1758 2290 1762
rect 2430 1758 2434 1762
rect 2694 1758 2698 1762
rect 3006 1758 3010 1762
rect 3086 1758 3090 1762
rect 158 1748 162 1752
rect 350 1748 354 1752
rect 398 1748 402 1752
rect 462 1748 466 1752
rect 662 1748 666 1752
rect 670 1748 674 1752
rect 686 1748 690 1752
rect 718 1748 722 1752
rect 750 1748 754 1752
rect 902 1748 906 1752
rect 1022 1748 1026 1752
rect 1262 1748 1266 1752
rect 1310 1748 1314 1752
rect 1366 1748 1370 1752
rect 1382 1748 1386 1752
rect 1398 1748 1402 1752
rect 1422 1748 1426 1752
rect 1478 1748 1482 1752
rect 1542 1748 1546 1752
rect 1830 1748 1834 1752
rect 1846 1748 1850 1752
rect 1862 1748 1866 1752
rect 1990 1748 1994 1752
rect 2150 1748 2154 1752
rect 2222 1748 2226 1752
rect 2254 1748 2258 1752
rect 2406 1748 2410 1752
rect 2462 1748 2466 1752
rect 2526 1748 2530 1752
rect 2574 1748 2578 1752
rect 2702 1748 2706 1752
rect 2814 1748 2818 1752
rect 2982 1748 2986 1752
rect 3070 1748 3074 1752
rect 3198 1748 3202 1752
rect 3438 1748 3442 1752
rect 3558 1748 3562 1752
rect 174 1738 178 1742
rect 230 1738 234 1742
rect 238 1738 242 1742
rect 494 1738 498 1742
rect 510 1738 514 1742
rect 542 1738 546 1742
rect 582 1738 586 1742
rect 606 1738 610 1742
rect 646 1738 650 1742
rect 654 1738 658 1742
rect 774 1738 778 1742
rect 1086 1738 1090 1742
rect 1110 1738 1114 1742
rect 1246 1738 1250 1742
rect 1422 1738 1426 1742
rect 1574 1738 1578 1742
rect 1710 1738 1714 1742
rect 1734 1738 1738 1742
rect 1822 1738 1826 1742
rect 1838 1738 1842 1742
rect 1926 1738 1930 1742
rect 2054 1738 2058 1742
rect 2134 1738 2138 1742
rect 2670 1738 2674 1742
rect 2806 1738 2810 1742
rect 3150 1738 3154 1742
rect 3406 1738 3410 1742
rect 3414 1738 3418 1742
rect 3494 1738 3498 1742
rect 3534 1738 3538 1742
rect 46 1728 50 1732
rect 238 1728 242 1732
rect 334 1728 338 1732
rect 926 1728 930 1732
rect 1038 1728 1042 1732
rect 1126 1728 1130 1732
rect 1206 1728 1210 1732
rect 1278 1728 1282 1732
rect 1390 1728 1394 1732
rect 1550 1728 1554 1732
rect 1574 1728 1578 1732
rect 1590 1728 1594 1732
rect 1606 1728 1610 1732
rect 1646 1728 1650 1732
rect 1710 1728 1714 1732
rect 1846 1728 1850 1732
rect 2022 1728 2026 1732
rect 2126 1728 2130 1732
rect 2134 1728 2138 1732
rect 2286 1728 2290 1732
rect 2310 1728 2314 1732
rect 2374 1728 2378 1732
rect 2422 1728 2426 1732
rect 3414 1728 3418 1732
rect 3502 1728 3506 1732
rect 102 1718 106 1722
rect 310 1718 314 1722
rect 318 1718 322 1722
rect 702 1718 706 1722
rect 1318 1718 1322 1722
rect 1358 1718 1362 1722
rect 1486 1718 1490 1722
rect 1654 1718 1658 1722
rect 1750 1718 1754 1722
rect 1766 1718 1770 1722
rect 1798 1718 1802 1722
rect 1822 1718 1826 1722
rect 1862 1718 1866 1722
rect 1870 1718 1874 1722
rect 2278 1718 2282 1722
rect 2574 1718 2578 1722
rect 2942 1718 2946 1722
rect 3478 1718 3482 1722
rect 3550 1718 3554 1722
rect 190 1708 194 1712
rect 238 1708 242 1712
rect 374 1708 378 1712
rect 558 1708 562 1712
rect 574 1708 578 1712
rect 590 1708 594 1712
rect 646 1708 650 1712
rect 726 1708 730 1712
rect 854 1708 858 1712
rect 1094 1708 1098 1712
rect 1126 1708 1130 1712
rect 1166 1708 1170 1712
rect 1198 1708 1202 1712
rect 1502 1708 1506 1712
rect 1742 1708 1746 1712
rect 1982 1708 1986 1712
rect 2118 1708 2122 1712
rect 2326 1708 2330 1712
rect 2350 1708 2354 1712
rect 2678 1708 2682 1712
rect 3030 1708 3034 1712
rect 3214 1708 3218 1712
rect 3526 1708 3530 1712
rect 994 1703 998 1707
rect 1002 1703 1005 1707
rect 1005 1703 1006 1707
rect 2026 1703 2030 1707
rect 2034 1703 2037 1707
rect 2037 1703 2038 1707
rect 3042 1703 3046 1707
rect 3050 1703 3053 1707
rect 3053 1703 3054 1707
rect 654 1698 658 1702
rect 1518 1698 1522 1702
rect 1790 1698 1794 1702
rect 1902 1698 1906 1702
rect 1998 1698 2002 1702
rect 2158 1698 2162 1702
rect 2350 1698 2354 1702
rect 2358 1698 2362 1702
rect 2510 1698 2514 1702
rect 2550 1698 2554 1702
rect 2614 1698 2618 1702
rect 2806 1698 2810 1702
rect 3470 1698 3474 1702
rect 278 1688 282 1692
rect 318 1688 322 1692
rect 350 1688 354 1692
rect 638 1688 642 1692
rect 782 1688 786 1692
rect 798 1688 802 1692
rect 814 1688 818 1692
rect 846 1688 850 1692
rect 966 1688 970 1692
rect 1038 1688 1042 1692
rect 1294 1688 1298 1692
rect 1302 1688 1306 1692
rect 1654 1688 1658 1692
rect 1718 1688 1722 1692
rect 1934 1688 1938 1692
rect 1950 1688 1954 1692
rect 1990 1688 1994 1692
rect 2086 1688 2090 1692
rect 2134 1688 2138 1692
rect 2238 1688 2242 1692
rect 2510 1688 2514 1692
rect 2542 1688 2546 1692
rect 2558 1688 2562 1692
rect 2590 1688 2594 1692
rect 694 1678 698 1682
rect 1062 1678 1066 1682
rect 1166 1678 1170 1682
rect 1198 1678 1202 1682
rect 2686 1688 2690 1692
rect 2974 1688 2978 1692
rect 3166 1688 3170 1692
rect 3182 1688 3186 1692
rect 3206 1688 3210 1692
rect 3254 1688 3258 1692
rect 3358 1688 3362 1692
rect 3366 1688 3370 1692
rect 3526 1688 3530 1692
rect 1742 1678 1746 1682
rect 1830 1678 1834 1682
rect 2006 1678 2010 1682
rect 2070 1678 2074 1682
rect 2102 1678 2106 1682
rect 2278 1678 2282 1682
rect 2318 1678 2322 1682
rect 2334 1678 2338 1682
rect 2350 1678 2354 1682
rect 2390 1678 2394 1682
rect 2406 1678 2410 1682
rect 2454 1678 2458 1682
rect 2710 1678 2714 1682
rect 2934 1678 2938 1682
rect 2974 1678 2978 1682
rect 3038 1678 3042 1682
rect 3350 1678 3354 1682
rect 3406 1678 3410 1682
rect 3518 1678 3522 1682
rect 3558 1678 3562 1682
rect 166 1668 170 1672
rect 294 1668 298 1672
rect 310 1668 314 1672
rect 422 1668 426 1672
rect 518 1668 522 1672
rect 678 1668 682 1672
rect 822 1668 826 1672
rect 1030 1668 1034 1672
rect 1054 1668 1058 1672
rect 1326 1668 1330 1672
rect 1342 1668 1346 1672
rect 1366 1668 1370 1672
rect 1406 1668 1410 1672
rect 1462 1668 1466 1672
rect 1518 1668 1522 1672
rect 1846 1668 1850 1672
rect 1934 1668 1938 1672
rect 1966 1668 1970 1672
rect 2110 1668 2114 1672
rect 2214 1668 2218 1672
rect 2270 1668 2274 1672
rect 2614 1668 2618 1672
rect 2902 1668 2906 1672
rect 3278 1668 3282 1672
rect 222 1658 226 1662
rect 254 1658 258 1662
rect 414 1658 418 1662
rect 582 1658 586 1662
rect 606 1658 610 1662
rect 622 1658 626 1662
rect 750 1658 754 1662
rect 766 1658 770 1662
rect 862 1658 866 1662
rect 870 1658 874 1662
rect 910 1658 914 1662
rect 1174 1658 1178 1662
rect 1182 1658 1186 1662
rect 1214 1658 1218 1662
rect 1278 1658 1282 1662
rect 1342 1658 1346 1662
rect 1414 1658 1418 1662
rect 1430 1658 1434 1662
rect 1454 1658 1458 1662
rect 1542 1658 1546 1662
rect 1606 1658 1610 1662
rect 1622 1658 1626 1662
rect 1678 1658 1682 1662
rect 1742 1658 1746 1662
rect 1766 1658 1770 1662
rect 1846 1658 1850 1662
rect 1878 1658 1882 1662
rect 1926 1658 1930 1662
rect 1958 1658 1962 1662
rect 1990 1658 1994 1662
rect 2174 1658 2178 1662
rect 2182 1658 2186 1662
rect 2190 1658 2194 1662
rect 2470 1658 2474 1662
rect 2526 1658 2530 1662
rect 2574 1658 2578 1662
rect 2630 1658 2634 1662
rect 2654 1658 2658 1662
rect 2774 1658 2778 1662
rect 2798 1658 2802 1662
rect 2878 1658 2882 1662
rect 3422 1658 3426 1662
rect 30 1648 34 1652
rect 158 1648 162 1652
rect 182 1648 186 1652
rect 422 1648 426 1652
rect 446 1648 450 1652
rect 486 1648 490 1652
rect 510 1648 514 1652
rect 774 1648 778 1652
rect 1254 1648 1258 1652
rect 1294 1648 1298 1652
rect 1430 1648 1434 1652
rect 1438 1648 1442 1652
rect 1582 1648 1586 1652
rect 1878 1648 1882 1652
rect 1910 1648 1914 1652
rect 1998 1648 2002 1652
rect 2102 1648 2106 1652
rect 2126 1648 2130 1652
rect 2206 1648 2210 1652
rect 2302 1648 2306 1652
rect 2422 1648 2426 1652
rect 2454 1648 2458 1652
rect 2662 1648 2666 1652
rect 2742 1648 2746 1652
rect 3182 1648 3186 1652
rect 3310 1648 3314 1652
rect 3326 1648 3330 1652
rect 3390 1648 3394 1652
rect 3470 1648 3474 1652
rect 342 1638 346 1642
rect 726 1638 730 1642
rect 1134 1638 1138 1642
rect 1254 1638 1258 1642
rect 2054 1638 2058 1642
rect 2110 1638 2114 1642
rect 2142 1638 2146 1642
rect 2238 1638 2242 1642
rect 2326 1638 2330 1642
rect 2598 1638 2602 1642
rect 2918 1638 2922 1642
rect 3294 1638 3298 1642
rect 158 1628 162 1632
rect 782 1628 786 1632
rect 1374 1628 1378 1632
rect 1382 1628 1386 1632
rect 1414 1628 1418 1632
rect 1614 1628 1618 1632
rect 1694 1628 1698 1632
rect 2270 1628 2274 1632
rect 2318 1628 2322 1632
rect 2334 1628 2338 1632
rect 2366 1628 2370 1632
rect 2422 1628 2426 1632
rect 2566 1628 2570 1632
rect 2886 1628 2890 1632
rect 398 1618 402 1622
rect 766 1618 770 1622
rect 1006 1618 1010 1622
rect 1126 1618 1130 1622
rect 238 1608 242 1612
rect 278 1608 282 1612
rect 438 1608 442 1612
rect 542 1608 546 1612
rect 1174 1618 1178 1622
rect 1358 1618 1362 1622
rect 1382 1618 1386 1622
rect 1598 1618 1602 1622
rect 1606 1618 1610 1622
rect 1726 1618 1730 1622
rect 1758 1618 1762 1622
rect 1870 1618 1874 1622
rect 2534 1618 2538 1622
rect 2638 1618 2642 1622
rect 2718 1618 2722 1622
rect 3134 1618 3138 1622
rect 886 1608 890 1612
rect 974 1608 978 1612
rect 1134 1608 1138 1612
rect 1150 1608 1154 1612
rect 1254 1608 1258 1612
rect 1262 1608 1266 1612
rect 1294 1608 1298 1612
rect 1398 1608 1402 1612
rect 1502 1608 1506 1612
rect 1638 1608 1642 1612
rect 1702 1608 1706 1612
rect 1734 1608 1738 1612
rect 1766 1608 1770 1612
rect 2686 1608 2690 1612
rect 2726 1608 2730 1612
rect 2758 1608 2762 1612
rect 3198 1608 3202 1612
rect 482 1603 486 1607
rect 490 1603 493 1607
rect 493 1603 494 1607
rect 1514 1603 1518 1607
rect 1522 1603 1525 1607
rect 1525 1603 1526 1607
rect 2538 1603 2542 1607
rect 2546 1603 2549 1607
rect 2549 1603 2550 1607
rect 190 1598 194 1602
rect 286 1598 290 1602
rect 310 1598 314 1602
rect 326 1598 330 1602
rect 390 1598 394 1602
rect 470 1598 474 1602
rect 638 1598 642 1602
rect 822 1598 826 1602
rect 1110 1598 1114 1602
rect 1350 1598 1354 1602
rect 1374 1598 1378 1602
rect 1550 1598 1554 1602
rect 1654 1598 1658 1602
rect 2486 1598 2490 1602
rect 2646 1598 2650 1602
rect 2710 1598 2714 1602
rect 2822 1598 2826 1602
rect 3326 1598 3330 1602
rect 534 1588 538 1592
rect 854 1588 858 1592
rect 1054 1588 1058 1592
rect 1294 1588 1298 1592
rect 1334 1588 1338 1592
rect 1366 1588 1370 1592
rect 1430 1588 1434 1592
rect 1478 1588 1482 1592
rect 2278 1588 2282 1592
rect 2358 1588 2362 1592
rect 2366 1588 2370 1592
rect 2462 1588 2466 1592
rect 2526 1588 2530 1592
rect 2862 1588 2866 1592
rect 2974 1588 2978 1592
rect 3062 1588 3066 1592
rect 3558 1588 3562 1592
rect 662 1578 666 1582
rect 710 1578 714 1582
rect 774 1578 778 1582
rect 926 1578 930 1582
rect 1102 1578 1106 1582
rect 1118 1578 1122 1582
rect 1286 1578 1290 1582
rect 1502 1578 1506 1582
rect 1574 1578 1578 1582
rect 1622 1578 1626 1582
rect 1638 1578 1642 1582
rect 1686 1578 1690 1582
rect 1710 1578 1714 1582
rect 1782 1578 1786 1582
rect 1798 1578 1802 1582
rect 2206 1578 2210 1582
rect 2222 1578 2226 1582
rect 2262 1578 2266 1582
rect 3462 1578 3466 1582
rect 206 1568 210 1572
rect 294 1568 298 1572
rect 326 1568 330 1572
rect 374 1568 378 1572
rect 414 1568 418 1572
rect 462 1568 466 1572
rect 534 1568 538 1572
rect 1142 1568 1146 1572
rect 1198 1568 1202 1572
rect 1230 1568 1234 1572
rect 1446 1568 1450 1572
rect 1494 1568 1498 1572
rect 1518 1568 1522 1572
rect 1590 1568 1594 1572
rect 1638 1568 1642 1572
rect 1702 1568 1706 1572
rect 1886 1568 1890 1572
rect 1894 1568 1898 1572
rect 2054 1568 2058 1572
rect 2142 1568 2146 1572
rect 2222 1568 2226 1572
rect 2238 1568 2242 1572
rect 2382 1568 2386 1572
rect 2502 1568 2506 1572
rect 2590 1568 2594 1572
rect 2742 1568 2746 1572
rect 2854 1568 2858 1572
rect 2942 1568 2946 1572
rect 3086 1568 3090 1572
rect 3158 1568 3162 1572
rect 3422 1568 3426 1572
rect 118 1558 122 1562
rect 150 1558 154 1562
rect 198 1558 202 1562
rect 374 1558 378 1562
rect 398 1558 402 1562
rect 718 1558 722 1562
rect 798 1558 802 1562
rect 886 1558 890 1562
rect 1054 1558 1058 1562
rect 1086 1558 1090 1562
rect 1342 1558 1346 1562
rect 1398 1558 1402 1562
rect 1430 1558 1434 1562
rect 1486 1558 1490 1562
rect 1534 1558 1538 1562
rect 1590 1558 1594 1562
rect 1606 1558 1610 1562
rect 1646 1558 1650 1562
rect 1742 1558 1746 1562
rect 1766 1558 1770 1562
rect 1830 1558 1834 1562
rect 1878 1558 1882 1562
rect 2038 1558 2042 1562
rect 2062 1558 2066 1562
rect 2294 1558 2298 1562
rect 2358 1558 2362 1562
rect 2422 1558 2426 1562
rect 2454 1558 2458 1562
rect 2582 1558 2586 1562
rect 2598 1558 2602 1562
rect 2662 1558 2666 1562
rect 2758 1558 2762 1562
rect 2894 1558 2898 1562
rect 2910 1558 2914 1562
rect 3070 1558 3074 1562
rect 3390 1558 3394 1562
rect 46 1548 50 1552
rect 222 1548 226 1552
rect 550 1548 554 1552
rect 582 1548 586 1552
rect 814 1548 818 1552
rect 1046 1548 1050 1552
rect 1222 1548 1226 1552
rect 1262 1548 1266 1552
rect 1470 1548 1474 1552
rect 1550 1548 1554 1552
rect 1574 1548 1578 1552
rect 1686 1548 1690 1552
rect 1694 1548 1698 1552
rect 1734 1548 1738 1552
rect 1846 1548 1850 1552
rect 1950 1548 1954 1552
rect 2046 1548 2050 1552
rect 2054 1548 2058 1552
rect 2134 1548 2138 1552
rect 2158 1548 2162 1552
rect 2262 1548 2266 1552
rect 2366 1548 2370 1552
rect 2390 1548 2394 1552
rect 2446 1548 2450 1552
rect 2550 1548 2554 1552
rect 2566 1548 2570 1552
rect 2598 1548 2602 1552
rect 2638 1548 2642 1552
rect 2846 1548 2850 1552
rect 2854 1548 2858 1552
rect 2870 1548 2874 1552
rect 2902 1548 2906 1552
rect 3062 1548 3066 1552
rect 3078 1548 3082 1552
rect 3534 1548 3538 1552
rect 3550 1548 3554 1552
rect 3558 1548 3562 1552
rect 286 1538 290 1542
rect 502 1538 506 1542
rect 526 1538 530 1542
rect 742 1538 746 1542
rect 870 1538 874 1542
rect 886 1538 890 1542
rect 942 1538 946 1542
rect 982 1538 986 1542
rect 1054 1538 1058 1542
rect 1334 1538 1338 1542
rect 1350 1538 1354 1542
rect 1414 1538 1418 1542
rect 1502 1538 1506 1542
rect 1606 1538 1610 1542
rect 1630 1538 1634 1542
rect 2094 1538 2098 1542
rect 2102 1538 2106 1542
rect 2150 1538 2154 1542
rect 2382 1538 2386 1542
rect 2398 1538 2402 1542
rect 2574 1538 2578 1542
rect 3470 1538 3474 1542
rect 150 1528 154 1532
rect 358 1528 362 1532
rect 366 1528 370 1532
rect 582 1528 586 1532
rect 614 1528 618 1532
rect 622 1528 626 1532
rect 910 1528 914 1532
rect 926 1528 930 1532
rect 1150 1528 1154 1532
rect 1182 1528 1186 1532
rect 1246 1528 1250 1532
rect 1342 1528 1346 1532
rect 1422 1528 1426 1532
rect 1478 1528 1482 1532
rect 1526 1528 1530 1532
rect 1550 1528 1554 1532
rect 1678 1528 1682 1532
rect 1806 1528 1810 1532
rect 1934 1528 1938 1532
rect 1982 1528 1986 1532
rect 2110 1528 2114 1532
rect 2222 1528 2226 1532
rect 2246 1528 2250 1532
rect 2262 1528 2266 1532
rect 2294 1528 2298 1532
rect 2342 1528 2346 1532
rect 2542 1528 2546 1532
rect 2646 1528 2650 1532
rect 2734 1528 2738 1532
rect 2758 1528 2762 1532
rect 2806 1528 2810 1532
rect 2814 1528 2818 1532
rect 2894 1528 2898 1532
rect 2926 1528 2930 1532
rect 2934 1528 2938 1532
rect 3142 1528 3146 1532
rect 3174 1528 3178 1532
rect 3342 1528 3346 1532
rect 174 1518 178 1522
rect 246 1518 250 1522
rect 398 1518 402 1522
rect 750 1518 754 1522
rect 1022 1518 1026 1522
rect 1150 1518 1154 1522
rect 1206 1518 1210 1522
rect 1262 1518 1266 1522
rect 1286 1518 1290 1522
rect 1382 1518 1386 1522
rect 1430 1518 1434 1522
rect 1462 1518 1466 1522
rect 1542 1518 1546 1522
rect 1558 1518 1562 1522
rect 1654 1518 1658 1522
rect 1686 1518 1690 1522
rect 1774 1518 1778 1522
rect 1822 1518 1826 1522
rect 1886 1518 1890 1522
rect 1910 1518 1914 1522
rect 1942 1518 1946 1522
rect 2006 1518 2010 1522
rect 2510 1518 2514 1522
rect 2574 1518 2578 1522
rect 2726 1518 2730 1522
rect 3182 1518 3186 1522
rect 3382 1518 3386 1522
rect 3430 1518 3434 1522
rect 110 1508 114 1512
rect 334 1508 338 1512
rect 630 1508 634 1512
rect 742 1508 746 1512
rect 862 1508 866 1512
rect 982 1508 986 1512
rect 1030 1508 1034 1512
rect 1166 1508 1170 1512
rect 1478 1508 1482 1512
rect 1646 1508 1650 1512
rect 1662 1508 1666 1512
rect 1694 1508 1698 1512
rect 1766 1508 1770 1512
rect 1838 1508 1842 1512
rect 1878 1508 1882 1512
rect 2014 1508 2018 1512
rect 2086 1508 2090 1512
rect 2150 1508 2154 1512
rect 2158 1508 2162 1512
rect 2854 1508 2858 1512
rect 2926 1508 2930 1512
rect 3126 1508 3130 1512
rect 3446 1508 3450 1512
rect 3462 1508 3466 1512
rect 994 1503 998 1507
rect 1002 1503 1005 1507
rect 1005 1503 1006 1507
rect 350 1498 354 1502
rect 358 1498 362 1502
rect 646 1498 650 1502
rect 766 1498 770 1502
rect 982 1498 986 1502
rect 1102 1498 1106 1502
rect 1246 1498 1250 1502
rect 1254 1498 1258 1502
rect 1270 1498 1274 1502
rect 1294 1498 1298 1502
rect 1350 1498 1354 1502
rect 1446 1498 1450 1502
rect 1614 1498 1618 1502
rect 1622 1498 1626 1502
rect 1646 1498 1650 1502
rect 2026 1503 2030 1507
rect 2034 1503 2037 1507
rect 2037 1503 2038 1507
rect 3042 1503 3046 1507
rect 3050 1503 3053 1507
rect 3053 1503 3054 1507
rect 1886 1498 1890 1502
rect 2094 1498 2098 1502
rect 2310 1498 2314 1502
rect 2478 1498 2482 1502
rect 2734 1498 2738 1502
rect 2790 1498 2794 1502
rect 2998 1498 3002 1502
rect 3230 1498 3234 1502
rect 438 1488 442 1492
rect 454 1488 458 1492
rect 822 1488 826 1492
rect 886 1488 890 1492
rect 1134 1488 1138 1492
rect 1198 1488 1202 1492
rect 1318 1488 1322 1492
rect 1414 1488 1418 1492
rect 1462 1488 1466 1492
rect 1638 1488 1642 1492
rect 1734 1488 1738 1492
rect 1758 1488 1762 1492
rect 1822 1488 1826 1492
rect 1838 1488 1842 1492
rect 2198 1488 2202 1492
rect 2286 1488 2290 1492
rect 2334 1488 2338 1492
rect 2358 1488 2362 1492
rect 2630 1488 2634 1492
rect 2662 1488 2666 1492
rect 3142 1488 3146 1492
rect 214 1478 218 1482
rect 414 1478 418 1482
rect 654 1478 658 1482
rect 838 1478 842 1482
rect 974 1478 978 1482
rect 1062 1478 1066 1482
rect 1166 1478 1170 1482
rect 1238 1478 1242 1482
rect 1334 1478 1338 1482
rect 1398 1478 1402 1482
rect 1414 1478 1418 1482
rect 1446 1478 1450 1482
rect 1454 1478 1458 1482
rect 1790 1478 1794 1482
rect 1814 1478 1818 1482
rect 1926 1478 1930 1482
rect 1990 1478 1994 1482
rect 2006 1478 2010 1482
rect 2134 1478 2138 1482
rect 2230 1478 2234 1482
rect 2270 1478 2274 1482
rect 2334 1478 2338 1482
rect 2366 1478 2370 1482
rect 2494 1478 2498 1482
rect 2878 1478 2882 1482
rect 2902 1478 2906 1482
rect 3294 1478 3298 1482
rect 3366 1478 3370 1482
rect 3422 1478 3426 1482
rect 3510 1478 3514 1482
rect 422 1468 426 1472
rect 814 1468 818 1472
rect 1022 1468 1026 1472
rect 1174 1468 1178 1472
rect 1238 1468 1242 1472
rect 1486 1468 1490 1472
rect 1510 1468 1514 1472
rect 1582 1468 1586 1472
rect 1606 1468 1610 1472
rect 1630 1468 1634 1472
rect 1766 1468 1770 1472
rect 1870 1468 1874 1472
rect 2182 1468 2186 1472
rect 2254 1468 2258 1472
rect 2358 1468 2362 1472
rect 2558 1468 2562 1472
rect 2582 1468 2586 1472
rect 2678 1468 2682 1472
rect 2742 1468 2746 1472
rect 2758 1468 2762 1472
rect 2894 1468 2898 1472
rect 2950 1468 2954 1472
rect 2982 1468 2986 1472
rect 3070 1468 3074 1472
rect 3334 1468 3338 1472
rect 3374 1468 3378 1472
rect 3406 1468 3410 1472
rect 3526 1468 3530 1472
rect 254 1458 258 1462
rect 262 1458 266 1462
rect 294 1458 298 1462
rect 694 1458 698 1462
rect 926 1458 930 1462
rect 966 1458 970 1462
rect 1054 1458 1058 1462
rect 1182 1458 1186 1462
rect 1262 1458 1266 1462
rect 1278 1458 1282 1462
rect 1302 1458 1306 1462
rect 1382 1458 1386 1462
rect 1446 1458 1450 1462
rect 1462 1458 1466 1462
rect 1534 1458 1538 1462
rect 1566 1458 1570 1462
rect 1622 1458 1626 1462
rect 1638 1458 1642 1462
rect 1726 1458 1730 1462
rect 1758 1458 1762 1462
rect 1902 1458 1906 1462
rect 2070 1458 2074 1462
rect 2142 1458 2146 1462
rect 2190 1458 2194 1462
rect 2198 1458 2202 1462
rect 2270 1458 2274 1462
rect 2278 1458 2282 1462
rect 2334 1458 2338 1462
rect 2550 1458 2554 1462
rect 2558 1458 2562 1462
rect 2686 1458 2690 1462
rect 2894 1458 2898 1462
rect 2926 1458 2930 1462
rect 3206 1458 3210 1462
rect 3246 1458 3250 1462
rect 3318 1458 3322 1462
rect 142 1448 146 1452
rect 158 1448 162 1452
rect 326 1448 330 1452
rect 606 1448 610 1452
rect 766 1448 770 1452
rect 830 1448 834 1452
rect 990 1448 994 1452
rect 1030 1448 1034 1452
rect 1086 1448 1090 1452
rect 1126 1448 1130 1452
rect 1270 1448 1274 1452
rect 1454 1448 1458 1452
rect 1542 1448 1546 1452
rect 1550 1448 1554 1452
rect 1590 1448 1594 1452
rect 1718 1448 1722 1452
rect 1750 1448 1754 1452
rect 1766 1448 1770 1452
rect 2030 1448 2034 1452
rect 2126 1448 2130 1452
rect 2206 1448 2210 1452
rect 2382 1448 2386 1452
rect 2422 1448 2426 1452
rect 2542 1448 2546 1452
rect 2566 1448 2570 1452
rect 2766 1448 2770 1452
rect 2886 1448 2890 1452
rect 2966 1448 2970 1452
rect 3214 1448 3218 1452
rect 3422 1448 3426 1452
rect 94 1438 98 1442
rect 390 1438 394 1442
rect 534 1438 538 1442
rect 822 1438 826 1442
rect 1006 1438 1010 1442
rect 1022 1438 1026 1442
rect 1062 1438 1066 1442
rect 1230 1438 1234 1442
rect 1286 1438 1290 1442
rect 1342 1438 1346 1442
rect 1414 1438 1418 1442
rect 1502 1438 1506 1442
rect 1726 1438 1730 1442
rect 1750 1438 1754 1442
rect 1934 1438 1938 1442
rect 2302 1438 2306 1442
rect 2366 1438 2370 1442
rect 2478 1438 2482 1442
rect 2790 1438 2794 1442
rect 3358 1438 3362 1442
rect 326 1428 330 1432
rect 446 1428 450 1432
rect 1006 1428 1010 1432
rect 1118 1428 1122 1432
rect 1774 1428 1778 1432
rect 2030 1428 2034 1432
rect 2078 1428 2082 1432
rect 2094 1428 2098 1432
rect 2238 1428 2242 1432
rect 310 1418 314 1422
rect 942 1418 946 1422
rect 1150 1418 1154 1422
rect 1206 1418 1210 1422
rect 1270 1418 1274 1422
rect 1294 1418 1298 1422
rect 1350 1418 1354 1422
rect 1422 1418 1426 1422
rect 1598 1418 1602 1422
rect 1694 1418 1698 1422
rect 1710 1418 1714 1422
rect 1742 1418 1746 1422
rect 1774 1418 1778 1422
rect 1846 1418 1850 1422
rect 2910 1418 2914 1422
rect 2990 1418 2994 1422
rect 3286 1418 3290 1422
rect 3358 1418 3362 1422
rect 318 1408 322 1412
rect 482 1403 486 1407
rect 490 1403 493 1407
rect 493 1403 494 1407
rect 1514 1403 1518 1407
rect 1522 1403 1525 1407
rect 1525 1403 1526 1407
rect 1942 1408 1946 1412
rect 2006 1408 2010 1412
rect 2102 1408 2106 1412
rect 2246 1408 2250 1412
rect 2406 1408 2410 1412
rect 2470 1408 2474 1412
rect 2590 1408 2594 1412
rect 2630 1408 2634 1412
rect 3430 1408 3434 1412
rect 2538 1403 2542 1407
rect 2546 1403 2549 1407
rect 2549 1403 2550 1407
rect 278 1398 282 1402
rect 558 1398 562 1402
rect 958 1398 962 1402
rect 998 1398 1002 1402
rect 1022 1398 1026 1402
rect 1302 1398 1306 1402
rect 1502 1398 1506 1402
rect 1582 1398 1586 1402
rect 1694 1398 1698 1402
rect 1718 1398 1722 1402
rect 1742 1398 1746 1402
rect 1806 1398 1810 1402
rect 1846 1398 1850 1402
rect 1870 1398 1874 1402
rect 1966 1398 1970 1402
rect 2054 1398 2058 1402
rect 2086 1398 2090 1402
rect 2166 1398 2170 1402
rect 2238 1398 2242 1402
rect 2446 1398 2450 1402
rect 2694 1398 2698 1402
rect 3390 1398 3394 1402
rect 246 1388 250 1392
rect 782 1388 786 1392
rect 870 1388 874 1392
rect 1078 1388 1082 1392
rect 1126 1388 1130 1392
rect 1158 1388 1162 1392
rect 1174 1388 1178 1392
rect 1246 1388 1250 1392
rect 1798 1388 1802 1392
rect 2078 1388 2082 1392
rect 2158 1388 2162 1392
rect 2166 1388 2170 1392
rect 2174 1388 2178 1392
rect 2190 1388 2194 1392
rect 2230 1388 2234 1392
rect 2294 1388 2298 1392
rect 2406 1388 2410 1392
rect 2574 1388 2578 1392
rect 2726 1388 2730 1392
rect 2862 1388 2866 1392
rect 3278 1388 3282 1392
rect 238 1378 242 1382
rect 358 1378 362 1382
rect 870 1378 874 1382
rect 910 1378 914 1382
rect 1022 1378 1026 1382
rect 1038 1378 1042 1382
rect 1086 1378 1090 1382
rect 1230 1378 1234 1382
rect 1638 1378 1642 1382
rect 1654 1378 1658 1382
rect 1822 1378 1826 1382
rect 1846 1378 1850 1382
rect 1910 1378 1914 1382
rect 2206 1378 2210 1382
rect 2350 1378 2354 1382
rect 2830 1378 2834 1382
rect 2902 1378 2906 1382
rect 3230 1378 3234 1382
rect 142 1368 146 1372
rect 166 1368 170 1372
rect 566 1368 570 1372
rect 942 1368 946 1372
rect 966 1368 970 1372
rect 1222 1368 1226 1372
rect 1662 1368 1666 1372
rect 1830 1368 1834 1372
rect 1894 1368 1898 1372
rect 1910 1368 1914 1372
rect 2030 1368 2034 1372
rect 2086 1368 2090 1372
rect 2142 1368 2146 1372
rect 2254 1368 2258 1372
rect 2390 1368 2394 1372
rect 2518 1368 2522 1372
rect 38 1358 42 1362
rect 310 1358 314 1362
rect 694 1358 698 1362
rect 1262 1358 1266 1362
rect 1342 1358 1346 1362
rect 1366 1358 1370 1362
rect 1494 1358 1498 1362
rect 1574 1358 1578 1362
rect 1606 1358 1610 1362
rect 1814 1358 1818 1362
rect 3134 1368 3138 1372
rect 1878 1358 1882 1362
rect 1918 1358 1922 1362
rect 2046 1358 2050 1362
rect 2190 1358 2194 1362
rect 2198 1358 2202 1362
rect 2366 1358 2370 1362
rect 2502 1358 2506 1362
rect 2526 1358 2530 1362
rect 2590 1358 2594 1362
rect 2686 1358 2690 1362
rect 2742 1358 2746 1362
rect 2758 1358 2762 1362
rect 3190 1358 3194 1362
rect 3334 1358 3338 1362
rect 446 1348 450 1352
rect 454 1348 458 1352
rect 502 1348 506 1352
rect 686 1348 690 1352
rect 846 1348 850 1352
rect 910 1348 914 1352
rect 1118 1348 1122 1352
rect 1182 1348 1186 1352
rect 1214 1348 1218 1352
rect 1342 1348 1346 1352
rect 1390 1348 1394 1352
rect 1398 1348 1402 1352
rect 1534 1348 1538 1352
rect 1582 1348 1586 1352
rect 1598 1348 1602 1352
rect 1630 1348 1634 1352
rect 1686 1348 1690 1352
rect 1766 1348 1770 1352
rect 1886 1348 1890 1352
rect 1942 1348 1946 1352
rect 1982 1348 1986 1352
rect 2054 1348 2058 1352
rect 2094 1348 2098 1352
rect 2214 1348 2218 1352
rect 2270 1348 2274 1352
rect 2398 1348 2402 1352
rect 2430 1348 2434 1352
rect 2502 1348 2506 1352
rect 2582 1348 2586 1352
rect 2614 1348 2618 1352
rect 2830 1348 2834 1352
rect 2854 1348 2858 1352
rect 2950 1348 2954 1352
rect 3006 1348 3010 1352
rect 3134 1348 3138 1352
rect 3454 1348 3458 1352
rect 342 1338 346 1342
rect 438 1338 442 1342
rect 942 1338 946 1342
rect 1006 1338 1010 1342
rect 1022 1338 1026 1342
rect 1086 1338 1090 1342
rect 1142 1338 1146 1342
rect 1326 1338 1330 1342
rect 1758 1338 1762 1342
rect 1830 1338 1834 1342
rect 1966 1338 1970 1342
rect 1990 1338 1994 1342
rect 2038 1338 2042 1342
rect 2270 1338 2274 1342
rect 2310 1338 2314 1342
rect 2510 1338 2514 1342
rect 2526 1338 2530 1342
rect 2582 1338 2586 1342
rect 2654 1338 2658 1342
rect 2702 1338 2706 1342
rect 2742 1338 2746 1342
rect 2758 1338 2762 1342
rect 2806 1338 2810 1342
rect 3110 1338 3114 1342
rect 3230 1338 3234 1342
rect 3270 1338 3274 1342
rect 3334 1338 3338 1342
rect 3358 1338 3362 1342
rect 3406 1338 3410 1342
rect 3430 1338 3434 1342
rect 358 1328 362 1332
rect 374 1328 378 1332
rect 742 1328 746 1332
rect 838 1328 842 1332
rect 950 1328 954 1332
rect 1030 1328 1034 1332
rect 1046 1328 1050 1332
rect 1150 1328 1154 1332
rect 1158 1328 1162 1332
rect 1206 1328 1210 1332
rect 1334 1328 1338 1332
rect 1366 1328 1370 1332
rect 1398 1328 1402 1332
rect 1406 1328 1410 1332
rect 1470 1328 1474 1332
rect 1566 1328 1570 1332
rect 1694 1328 1698 1332
rect 1734 1328 1738 1332
rect 1758 1328 1762 1332
rect 1846 1328 1850 1332
rect 1950 1328 1954 1332
rect 2102 1328 2106 1332
rect 2214 1328 2218 1332
rect 2222 1328 2226 1332
rect 2358 1328 2362 1332
rect 2366 1328 2370 1332
rect 2470 1328 2474 1332
rect 2598 1328 2602 1332
rect 2694 1328 2698 1332
rect 2766 1328 2770 1332
rect 2798 1328 2802 1332
rect 2918 1328 2922 1332
rect 2974 1328 2978 1332
rect 2998 1328 3002 1332
rect 3086 1328 3090 1332
rect 3302 1328 3306 1332
rect 3358 1328 3362 1332
rect 3422 1328 3426 1332
rect 3478 1328 3482 1332
rect 3502 1328 3506 1332
rect 350 1318 354 1322
rect 862 1318 866 1322
rect 1078 1318 1082 1322
rect 1342 1318 1346 1322
rect 1390 1318 1394 1322
rect 1414 1318 1418 1322
rect 1558 1318 1562 1322
rect 1694 1318 1698 1322
rect 1702 1318 1706 1322
rect 1822 1318 1826 1322
rect 1926 1318 1930 1322
rect 1934 1318 1938 1322
rect 2030 1318 2034 1322
rect 2046 1318 2050 1322
rect 2078 1318 2082 1322
rect 2118 1318 2122 1322
rect 2126 1318 2130 1322
rect 2166 1318 2170 1322
rect 2230 1318 2234 1322
rect 2246 1318 2250 1322
rect 2494 1318 2498 1322
rect 2510 1318 2514 1322
rect 2654 1318 2658 1322
rect 2702 1318 2706 1322
rect 2846 1318 2850 1322
rect 2926 1318 2930 1322
rect 3310 1318 3314 1322
rect 3350 1318 3354 1322
rect 526 1308 530 1312
rect 662 1308 666 1312
rect 846 1308 850 1312
rect 1102 1308 1106 1312
rect 1174 1308 1178 1312
rect 1606 1308 1610 1312
rect 1734 1308 1738 1312
rect 1782 1308 1786 1312
rect 1862 1308 1866 1312
rect 2094 1308 2098 1312
rect 2134 1308 2138 1312
rect 2350 1308 2354 1312
rect 2454 1308 2458 1312
rect 2470 1308 2474 1312
rect 2670 1308 2674 1312
rect 2990 1308 2994 1312
rect 3086 1308 3090 1312
rect 3358 1308 3362 1312
rect 994 1303 998 1307
rect 1002 1303 1005 1307
rect 1005 1303 1006 1307
rect 14 1298 18 1302
rect 406 1298 410 1302
rect 870 1298 874 1302
rect 1078 1298 1082 1302
rect 1142 1298 1146 1302
rect 1334 1298 1338 1302
rect 1382 1298 1386 1302
rect 1422 1298 1426 1302
rect 1582 1298 1586 1302
rect 1710 1298 1714 1302
rect 1750 1298 1754 1302
rect 1774 1298 1778 1302
rect 2026 1303 2030 1307
rect 2034 1303 2037 1307
rect 2037 1303 2038 1307
rect 1886 1298 1890 1302
rect 1902 1298 1906 1302
rect 2014 1298 2018 1302
rect 2182 1298 2186 1302
rect 2302 1298 2306 1302
rect 3042 1303 3046 1307
rect 3050 1303 3053 1307
rect 3053 1303 3054 1307
rect 2838 1298 2842 1302
rect 2854 1298 2858 1302
rect 2878 1298 2882 1302
rect 3030 1298 3034 1302
rect 3462 1298 3466 1302
rect 1030 1288 1034 1292
rect 1190 1288 1194 1292
rect 1254 1288 1258 1292
rect 1278 1288 1282 1292
rect 1294 1288 1298 1292
rect 1366 1288 1370 1292
rect 1398 1288 1402 1292
rect 1542 1288 1546 1292
rect 1558 1288 1562 1292
rect 1582 1288 1586 1292
rect 1598 1288 1602 1292
rect 1718 1288 1722 1292
rect 1798 1288 1802 1292
rect 1910 1288 1914 1292
rect 1974 1288 1978 1292
rect 2110 1288 2114 1292
rect 2174 1288 2178 1292
rect 2206 1288 2210 1292
rect 2246 1288 2250 1292
rect 2286 1288 2290 1292
rect 2454 1288 2458 1292
rect 2590 1288 2594 1292
rect 2614 1288 2618 1292
rect 3142 1288 3146 1292
rect 3318 1288 3322 1292
rect 3414 1288 3418 1292
rect 142 1278 146 1282
rect 166 1278 170 1282
rect 430 1278 434 1282
rect 622 1278 626 1282
rect 630 1278 634 1282
rect 854 1278 858 1282
rect 926 1278 930 1282
rect 1262 1278 1266 1282
rect 1278 1278 1282 1282
rect 1774 1278 1778 1282
rect 1822 1278 1826 1282
rect 1838 1278 1842 1282
rect 1862 1278 1866 1282
rect 2014 1278 2018 1282
rect 2118 1278 2122 1282
rect 2390 1278 2394 1282
rect 2406 1278 2410 1282
rect 2414 1278 2418 1282
rect 2926 1278 2930 1282
rect 2982 1278 2986 1282
rect 3190 1278 3194 1282
rect 3214 1278 3218 1282
rect 582 1268 586 1272
rect 614 1268 618 1272
rect 654 1268 658 1272
rect 750 1268 754 1272
rect 846 1268 850 1272
rect 870 1268 874 1272
rect 974 1268 978 1272
rect 1070 1268 1074 1272
rect 1078 1268 1082 1272
rect 1094 1268 1098 1272
rect 1286 1268 1290 1272
rect 1310 1268 1314 1272
rect 1358 1268 1362 1272
rect 1430 1268 1434 1272
rect 1462 1268 1466 1272
rect 1646 1268 1650 1272
rect 1670 1268 1674 1272
rect 1702 1268 1706 1272
rect 1758 1268 1762 1272
rect 1846 1268 1850 1272
rect 1894 1268 1898 1272
rect 1910 1268 1914 1272
rect 1934 1268 1938 1272
rect 1982 1268 1986 1272
rect 2022 1268 2026 1272
rect 2030 1268 2034 1272
rect 2094 1268 2098 1272
rect 2118 1268 2122 1272
rect 2142 1268 2146 1272
rect 2166 1268 2170 1272
rect 2246 1268 2250 1272
rect 2374 1268 2378 1272
rect 2390 1268 2394 1272
rect 2630 1268 2634 1272
rect 2638 1268 2642 1272
rect 2862 1268 2866 1272
rect 2878 1268 2882 1272
rect 2934 1268 2938 1272
rect 2974 1268 2978 1272
rect 3342 1268 3346 1272
rect 3486 1268 3490 1272
rect 102 1258 106 1262
rect 726 1258 730 1262
rect 782 1258 786 1262
rect 798 1258 802 1262
rect 814 1258 818 1262
rect 942 1258 946 1262
rect 982 1258 986 1262
rect 1030 1258 1034 1262
rect 1062 1258 1066 1262
rect 1102 1258 1106 1262
rect 1206 1258 1210 1262
rect 1318 1258 1322 1262
rect 1342 1258 1346 1262
rect 1374 1258 1378 1262
rect 1478 1258 1482 1262
rect 1550 1258 1554 1262
rect 1558 1258 1562 1262
rect 1574 1258 1578 1262
rect 1622 1258 1626 1262
rect 1638 1258 1642 1262
rect 1686 1258 1690 1262
rect 1710 1258 1714 1262
rect 1734 1258 1738 1262
rect 1742 1258 1746 1262
rect 1910 1258 1914 1262
rect 1942 1258 1946 1262
rect 2158 1258 2162 1262
rect 2446 1258 2450 1262
rect 2686 1258 2690 1262
rect 2718 1258 2722 1262
rect 2814 1258 2818 1262
rect 2926 1258 2930 1262
rect 2974 1258 2978 1262
rect 3422 1258 3426 1262
rect 198 1248 202 1252
rect 230 1248 234 1252
rect 238 1248 242 1252
rect 294 1248 298 1252
rect 310 1248 314 1252
rect 406 1248 410 1252
rect 654 1248 658 1252
rect 686 1248 690 1252
rect 766 1248 770 1252
rect 1086 1248 1090 1252
rect 1126 1248 1130 1252
rect 1222 1248 1226 1252
rect 1238 1248 1242 1252
rect 1318 1248 1322 1252
rect 1326 1248 1330 1252
rect 1366 1248 1370 1252
rect 1422 1248 1426 1252
rect 1806 1248 1810 1252
rect 1846 1248 1850 1252
rect 1854 1248 1858 1252
rect 2182 1248 2186 1252
rect 2342 1248 2346 1252
rect 2630 1248 2634 1252
rect 2710 1248 2714 1252
rect 2774 1248 2778 1252
rect 2838 1248 2842 1252
rect 3134 1248 3138 1252
rect 3278 1248 3282 1252
rect 374 1238 378 1242
rect 438 1238 442 1242
rect 926 1238 930 1242
rect 1078 1238 1082 1242
rect 1126 1238 1130 1242
rect 1278 1238 1282 1242
rect 1318 1238 1322 1242
rect 1614 1238 1618 1242
rect 1670 1238 1674 1242
rect 1766 1238 1770 1242
rect 1846 1238 1850 1242
rect 1990 1238 1994 1242
rect 2062 1238 2066 1242
rect 2078 1238 2082 1242
rect 2094 1238 2098 1242
rect 2198 1238 2202 1242
rect 2206 1238 2210 1242
rect 2270 1238 2274 1242
rect 2414 1238 2418 1242
rect 2430 1238 2434 1242
rect 2726 1238 2730 1242
rect 2742 1238 2746 1242
rect 2774 1238 2778 1242
rect 3070 1238 3074 1242
rect 638 1228 642 1232
rect 854 1228 858 1232
rect 1038 1228 1042 1232
rect 1054 1228 1058 1232
rect 1198 1228 1202 1232
rect 1206 1228 1210 1232
rect 1390 1228 1394 1232
rect 1414 1228 1418 1232
rect 1470 1228 1474 1232
rect 1550 1228 1554 1232
rect 1558 1228 1562 1232
rect 1654 1228 1658 1232
rect 1662 1228 1666 1232
rect 1774 1228 1778 1232
rect 1790 1228 1794 1232
rect 2142 1228 2146 1232
rect 2198 1228 2202 1232
rect 2286 1228 2290 1232
rect 2302 1228 2306 1232
rect 2806 1228 2810 1232
rect 646 1218 650 1222
rect 862 1218 866 1222
rect 1110 1218 1114 1222
rect 1286 1218 1290 1222
rect 1302 1218 1306 1222
rect 1342 1218 1346 1222
rect 1422 1218 1426 1222
rect 1894 1218 1898 1222
rect 1918 1218 1922 1222
rect 2046 1218 2050 1222
rect 2054 1218 2058 1222
rect 2422 1218 2426 1222
rect 1038 1208 1042 1212
rect 1430 1208 1434 1212
rect 1478 1208 1482 1212
rect 1870 1208 1874 1212
rect 1910 1208 1914 1212
rect 2014 1208 2018 1212
rect 2118 1208 2122 1212
rect 2334 1208 2338 1212
rect 2350 1208 2354 1212
rect 3126 1208 3130 1212
rect 482 1203 486 1207
rect 490 1203 493 1207
rect 493 1203 494 1207
rect 1514 1203 1518 1207
rect 1522 1203 1525 1207
rect 1525 1203 1526 1207
rect 2538 1203 2542 1207
rect 2546 1203 2549 1207
rect 2549 1203 2550 1207
rect 462 1198 466 1202
rect 726 1198 730 1202
rect 742 1198 746 1202
rect 958 1198 962 1202
rect 990 1198 994 1202
rect 1022 1198 1026 1202
rect 1070 1198 1074 1202
rect 1198 1198 1202 1202
rect 1254 1198 1258 1202
rect 1302 1198 1306 1202
rect 1334 1198 1338 1202
rect 2134 1198 2138 1202
rect 2638 1198 2642 1202
rect 2966 1198 2970 1202
rect 3182 1198 3186 1202
rect 3254 1198 3258 1202
rect 206 1188 210 1192
rect 390 1188 394 1192
rect 542 1188 546 1192
rect 942 1188 946 1192
rect 966 1188 970 1192
rect 1110 1188 1114 1192
rect 1318 1188 1322 1192
rect 1494 1188 1498 1192
rect 1598 1188 1602 1192
rect 1646 1188 1650 1192
rect 1710 1188 1714 1192
rect 1942 1188 1946 1192
rect 2030 1188 2034 1192
rect 2638 1188 2642 1192
rect 526 1178 530 1182
rect 1334 1178 1338 1182
rect 1390 1178 1394 1182
rect 1454 1178 1458 1182
rect 1750 1178 1754 1182
rect 1870 1178 1874 1182
rect 1918 1178 1922 1182
rect 1998 1178 2002 1182
rect 2086 1178 2090 1182
rect 2382 1178 2386 1182
rect 2646 1178 2650 1182
rect 942 1168 946 1172
rect 1238 1168 1242 1172
rect 1246 1168 1250 1172
rect 1270 1168 1274 1172
rect 1430 1168 1434 1172
rect 1462 1168 1466 1172
rect 1470 1168 1474 1172
rect 1494 1168 1498 1172
rect 1582 1168 1586 1172
rect 1718 1168 1722 1172
rect 1886 1168 1890 1172
rect 1926 1168 1930 1172
rect 2198 1168 2202 1172
rect 2622 1168 2626 1172
rect 2750 1168 2754 1172
rect 2758 1168 2762 1172
rect 2958 1168 2962 1172
rect 3094 1168 3098 1172
rect 3310 1168 3314 1172
rect 166 1158 170 1162
rect 286 1158 290 1162
rect 606 1158 610 1162
rect 678 1158 682 1162
rect 798 1158 802 1162
rect 822 1158 826 1162
rect 838 1158 842 1162
rect 1158 1158 1162 1162
rect 1318 1158 1322 1162
rect 1462 1158 1466 1162
rect 1510 1158 1514 1162
rect 1654 1158 1658 1162
rect 1670 1158 1674 1162
rect 1782 1158 1786 1162
rect 1806 1158 1810 1162
rect 1822 1158 1826 1162
rect 1862 1158 1866 1162
rect 1982 1158 1986 1162
rect 2062 1158 2066 1162
rect 2238 1158 2242 1162
rect 2310 1158 2314 1162
rect 2782 1158 2786 1162
rect 2982 1158 2986 1162
rect 3030 1158 3034 1162
rect 398 1148 402 1152
rect 518 1148 522 1152
rect 702 1148 706 1152
rect 718 1148 722 1152
rect 734 1148 738 1152
rect 750 1148 754 1152
rect 830 1148 834 1152
rect 998 1148 1002 1152
rect 1022 1148 1026 1152
rect 1086 1148 1090 1152
rect 1182 1148 1186 1152
rect 1222 1148 1226 1152
rect 1294 1148 1298 1152
rect 1302 1148 1306 1152
rect 1310 1148 1314 1152
rect 1478 1148 1482 1152
rect 1502 1148 1506 1152
rect 1534 1148 1538 1152
rect 1566 1148 1570 1152
rect 1686 1148 1690 1152
rect 1718 1148 1722 1152
rect 1774 1148 1778 1152
rect 1870 1148 1874 1152
rect 1886 1148 1890 1152
rect 1998 1148 2002 1152
rect 2022 1148 2026 1152
rect 2054 1148 2058 1152
rect 2142 1148 2146 1152
rect 2174 1148 2178 1152
rect 2254 1148 2258 1152
rect 2382 1148 2386 1152
rect 2614 1148 2618 1152
rect 3182 1148 3186 1152
rect 3558 1148 3562 1152
rect 6 1138 10 1142
rect 134 1138 138 1142
rect 838 1138 842 1142
rect 854 1138 858 1142
rect 862 1138 866 1142
rect 934 1138 938 1142
rect 1054 1138 1058 1142
rect 1230 1138 1234 1142
rect 1238 1138 1242 1142
rect 1550 1138 1554 1142
rect 1606 1138 1610 1142
rect 1614 1138 1618 1142
rect 1630 1138 1634 1142
rect 1654 1138 1658 1142
rect 1734 1138 1738 1142
rect 1854 1138 1858 1142
rect 1982 1138 1986 1142
rect 2070 1138 2074 1142
rect 2078 1138 2082 1142
rect 2478 1138 2482 1142
rect 2526 1138 2530 1142
rect 2702 1138 2706 1142
rect 2734 1138 2738 1142
rect 2846 1138 2850 1142
rect 2878 1138 2882 1142
rect 2958 1138 2962 1142
rect 3110 1138 3114 1142
rect 3302 1138 3306 1142
rect 3374 1138 3378 1142
rect 406 1128 410 1132
rect 462 1128 466 1132
rect 670 1128 674 1132
rect 742 1128 746 1132
rect 910 1128 914 1132
rect 926 1128 930 1132
rect 950 1128 954 1132
rect 1062 1128 1066 1132
rect 1302 1128 1306 1132
rect 1326 1128 1330 1132
rect 1334 1128 1338 1132
rect 1350 1128 1354 1132
rect 1430 1128 1434 1132
rect 1606 1128 1610 1132
rect 1646 1128 1650 1132
rect 1662 1128 1666 1132
rect 1798 1128 1802 1132
rect 1934 1128 1938 1132
rect 1942 1128 1946 1132
rect 2310 1128 2314 1132
rect 2478 1128 2482 1132
rect 2518 1128 2522 1132
rect 2542 1128 2546 1132
rect 2862 1128 2866 1132
rect 3030 1128 3034 1132
rect 3358 1128 3362 1132
rect 3382 1128 3386 1132
rect 766 1118 770 1122
rect 982 1118 986 1122
rect 1118 1118 1122 1122
rect 1182 1118 1186 1122
rect 1262 1118 1266 1122
rect 1342 1118 1346 1122
rect 1606 1118 1610 1122
rect 1622 1118 1626 1122
rect 1702 1118 1706 1122
rect 1814 1118 1818 1122
rect 1886 1118 1890 1122
rect 2070 1118 2074 1122
rect 2406 1118 2410 1122
rect 2662 1118 2666 1122
rect 3278 1118 3282 1122
rect 3302 1118 3306 1122
rect 3326 1118 3330 1122
rect 726 1108 730 1112
rect 822 1108 826 1112
rect 1110 1108 1114 1112
rect 1206 1108 1210 1112
rect 1222 1108 1226 1112
rect 1254 1108 1258 1112
rect 1286 1108 1290 1112
rect 1926 1108 1930 1112
rect 1958 1108 1962 1112
rect 1990 1108 1994 1112
rect 2110 1108 2114 1112
rect 2134 1108 2138 1112
rect 2774 1108 2778 1112
rect 3310 1108 3314 1112
rect 3494 1108 3498 1112
rect 994 1103 998 1107
rect 1002 1103 1005 1107
rect 1005 1103 1006 1107
rect 2026 1103 2030 1107
rect 2034 1103 2037 1107
rect 2037 1103 2038 1107
rect 3042 1103 3046 1107
rect 3050 1103 3053 1107
rect 3053 1103 3054 1107
rect 70 1098 74 1102
rect 390 1098 394 1102
rect 622 1098 626 1102
rect 654 1098 658 1102
rect 870 1098 874 1102
rect 910 1098 914 1102
rect 958 1098 962 1102
rect 1054 1098 1058 1102
rect 1174 1098 1178 1102
rect 1294 1098 1298 1102
rect 1406 1098 1410 1102
rect 1438 1098 1442 1102
rect 1486 1098 1490 1102
rect 1550 1098 1554 1102
rect 1638 1098 1642 1102
rect 1710 1098 1714 1102
rect 1726 1098 1730 1102
rect 1798 1098 1802 1102
rect 1806 1098 1810 1102
rect 1894 1098 1898 1102
rect 2046 1098 2050 1102
rect 2222 1098 2226 1102
rect 2262 1098 2266 1102
rect 2718 1098 2722 1102
rect 2774 1098 2778 1102
rect 2814 1098 2818 1102
rect 3062 1098 3066 1102
rect 3214 1098 3218 1102
rect 582 1088 586 1092
rect 774 1088 778 1092
rect 942 1088 946 1092
rect 990 1088 994 1092
rect 998 1088 1002 1092
rect 1030 1088 1034 1092
rect 1150 1088 1154 1092
rect 1190 1088 1194 1092
rect 1230 1088 1234 1092
rect 1310 1088 1314 1092
rect 1526 1088 1530 1092
rect 1534 1088 1538 1092
rect 1582 1088 1586 1092
rect 1590 1088 1594 1092
rect 1702 1088 1706 1092
rect 1830 1088 1834 1092
rect 2062 1088 2066 1092
rect 2150 1088 2154 1092
rect 2246 1088 2250 1092
rect 2262 1088 2266 1092
rect 2366 1088 2370 1092
rect 2398 1088 2402 1092
rect 2510 1088 2514 1092
rect 2998 1088 3002 1092
rect 3030 1088 3034 1092
rect 3278 1088 3282 1092
rect 86 1078 90 1082
rect 662 1078 666 1082
rect 886 1078 890 1082
rect 1126 1078 1130 1082
rect 1446 1078 1450 1082
rect 1462 1078 1466 1082
rect 1630 1078 1634 1082
rect 1734 1078 1738 1082
rect 1838 1078 1842 1082
rect 1934 1078 1938 1082
rect 2046 1078 2050 1082
rect 2070 1078 2074 1082
rect 2206 1078 2210 1082
rect 2214 1078 2218 1082
rect 2310 1078 2314 1082
rect 2558 1078 2562 1082
rect 2614 1078 2618 1082
rect 2726 1078 2730 1082
rect 2910 1078 2914 1082
rect 3222 1078 3226 1082
rect 358 1068 362 1072
rect 422 1068 426 1072
rect 566 1068 570 1072
rect 606 1068 610 1072
rect 798 1068 802 1072
rect 966 1068 970 1072
rect 974 1068 978 1072
rect 1022 1068 1026 1072
rect 1086 1068 1090 1072
rect 1134 1068 1138 1072
rect 1254 1068 1258 1072
rect 1262 1068 1266 1072
rect 1318 1068 1322 1072
rect 1374 1068 1378 1072
rect 1534 1068 1538 1072
rect 1590 1068 1594 1072
rect 1606 1068 1610 1072
rect 1662 1068 1666 1072
rect 1710 1068 1714 1072
rect 1766 1068 1770 1072
rect 1878 1068 1882 1072
rect 1950 1068 1954 1072
rect 1982 1068 1986 1072
rect 2006 1068 2010 1072
rect 2086 1068 2090 1072
rect 2110 1068 2114 1072
rect 2190 1068 2194 1072
rect 2230 1068 2234 1072
rect 2262 1068 2266 1072
rect 2414 1068 2418 1072
rect 2438 1068 2442 1072
rect 2550 1068 2554 1072
rect 2718 1068 2722 1072
rect 2926 1068 2930 1072
rect 2942 1068 2946 1072
rect 3182 1068 3186 1072
rect 222 1058 226 1062
rect 518 1058 522 1062
rect 622 1058 626 1062
rect 694 1058 698 1062
rect 710 1058 714 1062
rect 782 1058 786 1062
rect 830 1058 834 1062
rect 950 1058 954 1062
rect 1006 1058 1010 1062
rect 1030 1058 1034 1062
rect 1054 1058 1058 1062
rect 1070 1058 1074 1062
rect 1110 1058 1114 1062
rect 1126 1058 1130 1062
rect 1190 1058 1194 1062
rect 1214 1058 1218 1062
rect 1502 1058 1506 1062
rect 1526 1058 1530 1062
rect 1630 1058 1634 1062
rect 1894 1058 1898 1062
rect 1902 1058 1906 1062
rect 2094 1058 2098 1062
rect 2166 1058 2170 1062
rect 2326 1058 2330 1062
rect 2710 1058 2714 1062
rect 2918 1058 2922 1062
rect 3062 1058 3066 1062
rect 3382 1058 3386 1062
rect 22 1048 26 1052
rect 70 1048 74 1052
rect 822 1048 826 1052
rect 854 1048 858 1052
rect 886 1048 890 1052
rect 990 1048 994 1052
rect 1038 1048 1042 1052
rect 1054 1048 1058 1052
rect 1238 1048 1242 1052
rect 1398 1048 1402 1052
rect 1406 1048 1410 1052
rect 1510 1048 1514 1052
rect 1614 1048 1618 1052
rect 1646 1048 1650 1052
rect 1662 1048 1666 1052
rect 1694 1048 1698 1052
rect 1766 1048 1770 1052
rect 1902 1048 1906 1052
rect 1942 1048 1946 1052
rect 2062 1048 2066 1052
rect 2086 1048 2090 1052
rect 2254 1048 2258 1052
rect 2294 1048 2298 1052
rect 2302 1048 2306 1052
rect 2558 1048 2562 1052
rect 2854 1048 2858 1052
rect 3350 1048 3354 1052
rect 3374 1048 3378 1052
rect 6 1038 10 1042
rect 230 1038 234 1042
rect 438 1038 442 1042
rect 502 1038 506 1042
rect 574 1038 578 1042
rect 606 1038 610 1042
rect 654 1038 658 1042
rect 726 1038 730 1042
rect 1174 1038 1178 1042
rect 1294 1038 1298 1042
rect 1326 1038 1330 1042
rect 1350 1038 1354 1042
rect 1526 1038 1530 1042
rect 1686 1038 1690 1042
rect 1966 1038 1970 1042
rect 2222 1038 2226 1042
rect 2494 1038 2498 1042
rect 3214 1038 3218 1042
rect 3430 1038 3434 1042
rect 206 1028 210 1032
rect 590 1028 594 1032
rect 910 1028 914 1032
rect 934 1028 938 1032
rect 974 1028 978 1032
rect 1094 1028 1098 1032
rect 1406 1028 1410 1032
rect 1422 1028 1426 1032
rect 1462 1028 1466 1032
rect 1558 1028 1562 1032
rect 2150 1028 2154 1032
rect 2518 1028 2522 1032
rect 2918 1028 2922 1032
rect 3366 1028 3370 1032
rect 3470 1028 3474 1032
rect 134 1018 138 1022
rect 1094 1018 1098 1022
rect 1102 1018 1106 1022
rect 1174 1018 1178 1022
rect 1182 1018 1186 1022
rect 1446 1018 1450 1022
rect 1494 1018 1498 1022
rect 1670 1018 1674 1022
rect 1990 1018 1994 1022
rect 2022 1018 2026 1022
rect 2974 1018 2978 1022
rect 3054 1018 3058 1022
rect 862 1008 866 1012
rect 1062 1008 1066 1012
rect 1334 1008 1338 1012
rect 1390 1008 1394 1012
rect 1398 1008 1402 1012
rect 1486 1008 1490 1012
rect 1494 1008 1498 1012
rect 1598 1008 1602 1012
rect 1894 1008 1898 1012
rect 2118 1008 2122 1012
rect 2270 1008 2274 1012
rect 2286 1008 2290 1012
rect 2294 1008 2298 1012
rect 2342 1008 2346 1012
rect 2958 1008 2962 1012
rect 482 1003 486 1007
rect 490 1003 493 1007
rect 493 1003 494 1007
rect 1514 1003 1518 1007
rect 1522 1003 1525 1007
rect 1525 1003 1526 1007
rect 2538 1003 2542 1007
rect 2546 1003 2549 1007
rect 2549 1003 2550 1007
rect 782 998 786 1002
rect 974 998 978 1002
rect 1062 998 1066 1002
rect 1086 998 1090 1002
rect 1182 998 1186 1002
rect 1326 998 1330 1002
rect 1470 998 1474 1002
rect 1598 998 1602 1002
rect 1686 998 1690 1002
rect 1734 998 1738 1002
rect 2062 998 2066 1002
rect 2206 998 2210 1002
rect 2486 998 2490 1002
rect 3510 998 3514 1002
rect 366 988 370 992
rect 534 988 538 992
rect 734 988 738 992
rect 870 988 874 992
rect 998 988 1002 992
rect 1006 988 1010 992
rect 1206 988 1210 992
rect 1246 988 1250 992
rect 1358 988 1362 992
rect 1910 988 1914 992
rect 1982 988 1986 992
rect 2238 988 2242 992
rect 2422 988 2426 992
rect 3526 988 3530 992
rect 470 978 474 982
rect 510 978 514 982
rect 742 978 746 982
rect 1174 978 1178 982
rect 1454 978 1458 982
rect 1478 978 1482 982
rect 1918 978 1922 982
rect 2598 978 2602 982
rect 2606 978 2610 982
rect 2926 978 2930 982
rect 2966 978 2970 982
rect 3238 978 3242 982
rect 3510 978 3514 982
rect 1054 968 1058 972
rect 1118 968 1122 972
rect 1150 968 1154 972
rect 1182 968 1186 972
rect 1230 968 1234 972
rect 1398 968 1402 972
rect 1406 968 1410 972
rect 1558 968 1562 972
rect 1590 968 1594 972
rect 1646 968 1650 972
rect 1670 968 1674 972
rect 1870 968 1874 972
rect 1950 968 1954 972
rect 1958 968 1962 972
rect 2110 968 2114 972
rect 2190 968 2194 972
rect 2238 968 2242 972
rect 2262 968 2266 972
rect 2350 968 2354 972
rect 2894 968 2898 972
rect 3342 968 3346 972
rect 3374 968 3378 972
rect 3542 968 3546 972
rect 6 958 10 962
rect 86 958 90 962
rect 294 958 298 962
rect 382 958 386 962
rect 630 958 634 962
rect 694 958 698 962
rect 790 958 794 962
rect 830 958 834 962
rect 1102 958 1106 962
rect 1126 958 1130 962
rect 1142 958 1146 962
rect 1262 958 1266 962
rect 1398 958 1402 962
rect 1758 958 1762 962
rect 1798 958 1802 962
rect 1998 958 2002 962
rect 2014 958 2018 962
rect 2182 958 2186 962
rect 2206 958 2210 962
rect 2766 958 2770 962
rect 3086 958 3090 962
rect 3470 958 3474 962
rect 414 948 418 952
rect 646 948 650 952
rect 678 948 682 952
rect 910 948 914 952
rect 1006 948 1010 952
rect 1046 948 1050 952
rect 1134 948 1138 952
rect 1150 948 1154 952
rect 1214 948 1218 952
rect 1222 948 1226 952
rect 1262 948 1266 952
rect 1334 948 1338 952
rect 1510 948 1514 952
rect 1574 948 1578 952
rect 1582 948 1586 952
rect 1662 948 1666 952
rect 1870 948 1874 952
rect 1902 948 1906 952
rect 1966 948 1970 952
rect 2030 948 2034 952
rect 2158 948 2162 952
rect 2182 948 2186 952
rect 2366 948 2370 952
rect 2390 948 2394 952
rect 2654 948 2658 952
rect 2982 948 2986 952
rect 3094 948 3098 952
rect 3214 948 3218 952
rect 3230 948 3234 952
rect 3382 948 3386 952
rect 3422 948 3426 952
rect 182 938 186 942
rect 254 938 258 942
rect 318 938 322 942
rect 470 938 474 942
rect 614 938 618 942
rect 774 938 778 942
rect 846 938 850 942
rect 862 938 866 942
rect 870 938 874 942
rect 910 938 914 942
rect 982 938 986 942
rect 1038 938 1042 942
rect 1054 938 1058 942
rect 1198 938 1202 942
rect 1254 938 1258 942
rect 1422 938 1426 942
rect 1454 938 1458 942
rect 1678 938 1682 942
rect 1686 938 1690 942
rect 1782 938 1786 942
rect 1798 938 1802 942
rect 1806 938 1810 942
rect 1846 940 1850 942
rect 1846 938 1850 940
rect 1854 938 1858 942
rect 2062 938 2066 942
rect 2166 938 2170 942
rect 2198 938 2202 942
rect 2326 938 2330 942
rect 2374 938 2378 942
rect 3238 938 3242 942
rect 3270 938 3274 942
rect 278 928 282 932
rect 782 928 786 932
rect 942 928 946 932
rect 1094 928 1098 932
rect 1182 928 1186 932
rect 1238 928 1242 932
rect 1278 928 1282 932
rect 1302 928 1306 932
rect 1350 928 1354 932
rect 1374 928 1378 932
rect 1414 928 1418 932
rect 1590 928 1594 932
rect 1670 928 1674 932
rect 1726 928 1730 932
rect 1822 928 1826 932
rect 1838 928 1842 932
rect 2046 928 2050 932
rect 2086 928 2090 932
rect 2390 928 2394 932
rect 3054 928 3058 932
rect 3070 928 3074 932
rect 3222 928 3226 932
rect 230 918 234 922
rect 630 918 634 922
rect 726 918 730 922
rect 774 918 778 922
rect 926 918 930 922
rect 982 918 986 922
rect 1038 918 1042 922
rect 1166 918 1170 922
rect 1342 918 1346 922
rect 1550 918 1554 922
rect 1710 918 1714 922
rect 1750 918 1754 922
rect 1950 918 1954 922
rect 1974 918 1978 922
rect 2062 918 2066 922
rect 2102 918 2106 922
rect 2310 918 2314 922
rect 2710 918 2714 922
rect 254 908 258 912
rect 542 908 546 912
rect 1078 908 1082 912
rect 1238 908 1242 912
rect 1254 908 1258 912
rect 1302 908 1306 912
rect 1438 908 1442 912
rect 1702 908 1706 912
rect 1798 908 1802 912
rect 1894 908 1898 912
rect 1918 908 1922 912
rect 1934 908 1938 912
rect 2230 908 2234 912
rect 2638 908 2642 912
rect 2718 908 2722 912
rect 2894 908 2898 912
rect 3102 908 3106 912
rect 994 903 998 907
rect 1002 903 1005 907
rect 1005 903 1006 907
rect 2026 903 2030 907
rect 2034 903 2037 907
rect 2037 903 2038 907
rect 782 898 786 902
rect 790 898 794 902
rect 862 898 866 902
rect 982 898 986 902
rect 1030 898 1034 902
rect 1214 898 1218 902
rect 2134 898 2138 902
rect 2350 898 2354 902
rect 3042 903 3046 907
rect 3050 903 3053 907
rect 3053 903 3054 907
rect 462 888 466 892
rect 790 888 794 892
rect 854 888 858 892
rect 990 888 994 892
rect 1110 888 1114 892
rect 1174 888 1178 892
rect 1206 888 1210 892
rect 1238 888 1242 892
rect 1254 888 1258 892
rect 1470 888 1474 892
rect 1558 888 1562 892
rect 1742 888 1746 892
rect 1750 888 1754 892
rect 1942 888 1946 892
rect 1958 888 1962 892
rect 1982 888 1986 892
rect 2046 888 2050 892
rect 2102 888 2106 892
rect 2262 888 2266 892
rect 2278 888 2282 892
rect 2614 888 2618 892
rect 2966 888 2970 892
rect 3030 888 3034 892
rect 3046 888 3050 892
rect 54 878 58 882
rect 622 878 626 882
rect 798 878 802 882
rect 998 878 1002 882
rect 1022 878 1026 882
rect 1150 878 1154 882
rect 1158 878 1162 882
rect 1270 878 1274 882
rect 1278 878 1282 882
rect 1478 878 1482 882
rect 1694 878 1698 882
rect 2310 878 2314 882
rect 2462 878 2466 882
rect 2854 878 2858 882
rect 2982 878 2986 882
rect 558 868 562 872
rect 686 868 690 872
rect 694 868 698 872
rect 902 868 906 872
rect 990 868 994 872
rect 1030 868 1034 872
rect 1174 868 1178 872
rect 1182 868 1186 872
rect 1230 868 1234 872
rect 1310 868 1314 872
rect 1334 868 1338 872
rect 1422 868 1426 872
rect 1486 868 1490 872
rect 1606 868 1610 872
rect 1702 868 1706 872
rect 1814 868 1818 872
rect 2038 868 2042 872
rect 2054 868 2058 872
rect 2118 868 2122 872
rect 2150 868 2154 872
rect 2198 868 2202 872
rect 2246 868 2250 872
rect 2302 868 2306 872
rect 2446 868 2450 872
rect 2510 868 2514 872
rect 2518 868 2522 872
rect 238 858 242 862
rect 286 858 290 862
rect 334 858 338 862
rect 350 858 354 862
rect 446 858 450 862
rect 614 858 618 862
rect 622 858 626 862
rect 718 858 722 862
rect 758 858 762 862
rect 806 858 810 862
rect 838 858 842 862
rect 862 858 866 862
rect 870 858 874 862
rect 950 858 954 862
rect 1142 858 1146 862
rect 1318 858 1322 862
rect 1342 858 1346 862
rect 1390 858 1394 862
rect 1398 858 1402 862
rect 1558 858 1562 862
rect 1566 858 1570 862
rect 1590 858 1594 862
rect 1670 858 1674 862
rect 1726 858 1730 862
rect 1942 858 1946 862
rect 2406 858 2410 862
rect 2430 858 2434 862
rect 2686 858 2690 862
rect 2870 858 2874 862
rect 2902 858 2906 862
rect 286 848 290 852
rect 582 848 586 852
rect 670 848 674 852
rect 878 848 882 852
rect 966 848 970 852
rect 982 848 986 852
rect 1110 848 1114 852
rect 1118 848 1122 852
rect 1174 848 1178 852
rect 1206 848 1210 852
rect 1294 848 1298 852
rect 1390 848 1394 852
rect 1414 848 1418 852
rect 1430 848 1434 852
rect 1462 848 1466 852
rect 1470 848 1474 852
rect 1550 848 1554 852
rect 1574 848 1578 852
rect 1670 848 1674 852
rect 1822 848 1826 852
rect 1926 848 1930 852
rect 1958 848 1962 852
rect 2046 848 2050 852
rect 2086 848 2090 852
rect 2238 848 2242 852
rect 3102 848 3106 852
rect 3222 848 3226 852
rect 118 838 122 842
rect 446 838 450 842
rect 518 838 522 842
rect 590 838 594 842
rect 702 838 706 842
rect 718 838 722 842
rect 974 838 978 842
rect 1054 838 1058 842
rect 1302 838 1306 842
rect 1374 838 1378 842
rect 1438 838 1442 842
rect 1446 838 1450 842
rect 1478 838 1482 842
rect 1910 838 1914 842
rect 2070 838 2074 842
rect 2158 838 2162 842
rect 2294 838 2298 842
rect 2670 838 2674 842
rect 2710 838 2714 842
rect 3118 838 3122 842
rect 3166 838 3170 842
rect 62 828 66 832
rect 606 828 610 832
rect 1054 828 1058 832
rect 1110 828 1114 832
rect 1238 828 1242 832
rect 1550 828 1554 832
rect 1558 828 1562 832
rect 1574 828 1578 832
rect 1606 828 1610 832
rect 566 818 570 822
rect 1894 818 1898 822
rect 2022 818 2026 822
rect 2038 818 2042 822
rect 2286 818 2290 822
rect 2446 818 2450 822
rect 2678 818 2682 822
rect 2702 818 2706 822
rect 206 808 210 812
rect 334 808 338 812
rect 350 808 354 812
rect 462 808 466 812
rect 974 808 978 812
rect 990 808 994 812
rect 1262 808 1266 812
rect 1382 808 1386 812
rect 1390 808 1394 812
rect 1758 808 1762 812
rect 3094 808 3098 812
rect 482 803 486 807
rect 490 803 493 807
rect 493 803 494 807
rect 1514 803 1518 807
rect 1522 803 1525 807
rect 1525 803 1526 807
rect 2538 803 2542 807
rect 2546 803 2549 807
rect 2549 803 2550 807
rect 182 798 186 802
rect 454 798 458 802
rect 590 798 594 802
rect 766 798 770 802
rect 790 798 794 802
rect 1246 798 1250 802
rect 1254 798 1258 802
rect 1310 798 1314 802
rect 1494 798 1498 802
rect 1638 798 1642 802
rect 1798 798 1802 802
rect 2390 798 2394 802
rect 2526 798 2530 802
rect 2566 798 2570 802
rect 734 788 738 792
rect 990 788 994 792
rect 1166 788 1170 792
rect 1198 788 1202 792
rect 1334 788 1338 792
rect 1350 788 1354 792
rect 1374 788 1378 792
rect 1390 788 1394 792
rect 1510 788 1514 792
rect 1542 788 1546 792
rect 1670 788 1674 792
rect 1710 788 1714 792
rect 1902 788 1906 792
rect 2438 788 2442 792
rect 2598 788 2602 792
rect 822 778 826 782
rect 830 778 834 782
rect 1158 778 1162 782
rect 1342 778 1346 782
rect 2566 778 2570 782
rect 2630 778 2634 782
rect 2902 778 2906 782
rect 3462 778 3466 782
rect 462 768 466 772
rect 1134 768 1138 772
rect 1206 768 1210 772
rect 1574 768 1578 772
rect 1614 768 1618 772
rect 1638 768 1642 772
rect 1774 768 1778 772
rect 2046 768 2050 772
rect 2054 768 2058 772
rect 2094 768 2098 772
rect 2110 768 2114 772
rect 2734 768 2738 772
rect 3534 768 3538 772
rect 302 758 306 762
rect 710 758 714 762
rect 718 758 722 762
rect 838 758 842 762
rect 998 758 1002 762
rect 1070 758 1074 762
rect 1142 758 1146 762
rect 1230 758 1234 762
rect 1238 758 1242 762
rect 1286 758 1290 762
rect 1350 758 1354 762
rect 1598 758 1602 762
rect 1830 758 1834 762
rect 1982 758 1986 762
rect 2158 758 2162 762
rect 2334 758 2338 762
rect 2406 758 2410 762
rect 3094 758 3098 762
rect 3166 758 3170 762
rect 582 748 586 752
rect 606 748 610 752
rect 726 748 730 752
rect 854 748 858 752
rect 1590 748 1594 752
rect 1622 748 1626 752
rect 1726 748 1730 752
rect 1838 748 1842 752
rect 1862 748 1866 752
rect 1998 748 2002 752
rect 2134 748 2138 752
rect 2174 748 2178 752
rect 2198 748 2202 752
rect 2286 748 2290 752
rect 2758 748 2762 752
rect 2838 748 2842 752
rect 182 738 186 742
rect 318 738 322 742
rect 510 738 514 742
rect 574 738 578 742
rect 766 738 770 742
rect 814 738 818 742
rect 878 738 882 742
rect 1198 738 1202 742
rect 1286 738 1290 742
rect 1310 738 1314 742
rect 1326 738 1330 742
rect 1342 738 1346 742
rect 1406 738 1410 742
rect 1414 738 1418 742
rect 1430 738 1434 742
rect 1654 738 1658 742
rect 1726 738 1730 742
rect 1734 738 1738 742
rect 1782 738 1786 742
rect 1830 738 1834 742
rect 1958 738 1962 742
rect 2006 738 2010 742
rect 2022 738 2026 742
rect 2230 738 2234 742
rect 2270 738 2274 742
rect 2470 738 2474 742
rect 2902 748 2906 752
rect 2726 738 2730 742
rect 2750 738 2754 742
rect 2766 738 2770 742
rect 2974 738 2978 742
rect 2998 738 3002 742
rect 3078 738 3082 742
rect 3094 738 3098 742
rect 3294 738 3298 742
rect 374 728 378 732
rect 558 728 562 732
rect 582 728 586 732
rect 710 728 714 732
rect 886 728 890 732
rect 950 728 954 732
rect 974 728 978 732
rect 1030 728 1034 732
rect 1230 728 1234 732
rect 1238 728 1242 732
rect 1582 728 1586 732
rect 1782 728 1786 732
rect 1950 728 1954 732
rect 2054 728 2058 732
rect 2118 728 2122 732
rect 2318 728 2322 732
rect 2414 728 2418 732
rect 2478 728 2482 732
rect 2622 728 2626 732
rect 2654 728 2658 732
rect 2958 728 2962 732
rect 3038 728 3042 732
rect 3222 728 3226 732
rect 414 718 418 722
rect 542 718 546 722
rect 558 718 562 722
rect 654 718 658 722
rect 1454 718 1458 722
rect 1486 718 1490 722
rect 1494 718 1498 722
rect 1566 718 1570 722
rect 1590 718 1594 722
rect 1622 718 1626 722
rect 1854 718 1858 722
rect 1934 718 1938 722
rect 2158 718 2162 722
rect 2286 718 2290 722
rect 2366 718 2370 722
rect 2870 718 2874 722
rect 38 708 42 712
rect 182 708 186 712
rect 262 708 266 712
rect 438 708 442 712
rect 878 708 882 712
rect 886 708 890 712
rect 1110 708 1114 712
rect 1158 708 1162 712
rect 1174 708 1178 712
rect 1286 708 1290 712
rect 1446 708 1450 712
rect 1478 708 1482 712
rect 1558 708 1562 712
rect 1646 708 1650 712
rect 2014 708 2018 712
rect 2342 708 2346 712
rect 2566 708 2570 712
rect 2886 708 2890 712
rect 994 703 998 707
rect 1002 703 1005 707
rect 1005 703 1006 707
rect 2026 703 2030 707
rect 2034 703 2037 707
rect 2037 703 2038 707
rect 3042 703 3046 707
rect 3050 703 3053 707
rect 3053 703 3054 707
rect 158 698 162 702
rect 246 698 250 702
rect 590 698 594 702
rect 726 698 730 702
rect 742 698 746 702
rect 982 698 986 702
rect 1038 698 1042 702
rect 1238 698 1242 702
rect 1798 698 1802 702
rect 2014 698 2018 702
rect 2174 698 2178 702
rect 2390 698 2394 702
rect 2910 698 2914 702
rect 3222 698 3226 702
rect 310 688 314 692
rect 718 688 722 692
rect 774 688 778 692
rect 910 688 914 692
rect 1206 688 1210 692
rect 1318 688 1322 692
rect 1582 688 1586 692
rect 1710 688 1714 692
rect 1734 688 1738 692
rect 1758 688 1762 692
rect 1814 688 1818 692
rect 1830 688 1834 692
rect 1870 688 1874 692
rect 2318 688 2322 692
rect 2398 688 2402 692
rect 2598 688 2602 692
rect 2990 688 2994 692
rect 3150 688 3154 692
rect 3206 688 3210 692
rect 3214 688 3218 692
rect 470 678 474 682
rect 518 678 522 682
rect 726 678 730 682
rect 966 678 970 682
rect 1070 678 1074 682
rect 1086 678 1090 682
rect 1126 678 1130 682
rect 1134 678 1138 682
rect 1150 678 1154 682
rect 1230 678 1234 682
rect 1278 678 1282 682
rect 1326 678 1330 682
rect 1342 678 1346 682
rect 1358 678 1362 682
rect 1398 678 1402 682
rect 1430 678 1434 682
rect 1502 678 1506 682
rect 1518 678 1522 682
rect 1614 678 1618 682
rect 1654 678 1658 682
rect 1726 678 1730 682
rect 1910 678 1914 682
rect 2014 678 2018 682
rect 2070 678 2074 682
rect 2126 678 2130 682
rect 2310 678 2314 682
rect 2406 678 2410 682
rect 2526 678 2530 682
rect 3102 678 3106 682
rect 3222 678 3226 682
rect 126 668 130 672
rect 374 668 378 672
rect 670 668 674 672
rect 686 668 690 672
rect 734 668 738 672
rect 838 668 842 672
rect 1030 668 1034 672
rect 1510 668 1514 672
rect 1702 668 1706 672
rect 1782 668 1786 672
rect 1790 668 1794 672
rect 1886 668 1890 672
rect 2110 668 2114 672
rect 2206 668 2210 672
rect 2374 668 2378 672
rect 2430 668 2434 672
rect 2438 668 2442 672
rect 3062 668 3066 672
rect 3214 668 3218 672
rect 302 658 306 662
rect 334 658 338 662
rect 382 658 386 662
rect 446 658 450 662
rect 470 658 474 662
rect 526 658 530 662
rect 750 658 754 662
rect 790 658 794 662
rect 958 658 962 662
rect 1238 658 1242 662
rect 1246 658 1250 662
rect 1278 658 1282 662
rect 1286 658 1290 662
rect 1398 658 1402 662
rect 1758 658 1762 662
rect 1766 658 1770 662
rect 1854 658 1858 662
rect 1886 658 1890 662
rect 1926 658 1930 662
rect 2062 658 2066 662
rect 2086 658 2090 662
rect 2134 658 2138 662
rect 2150 658 2154 662
rect 2342 658 2346 662
rect 2646 658 2650 662
rect 2742 658 2746 662
rect 2790 658 2794 662
rect 2886 658 2890 662
rect 3246 658 3250 662
rect 198 648 202 652
rect 382 648 386 652
rect 390 648 394 652
rect 518 648 522 652
rect 590 648 594 652
rect 654 648 658 652
rect 710 648 714 652
rect 726 648 730 652
rect 1366 648 1370 652
rect 1454 648 1458 652
rect 1542 648 1546 652
rect 1550 648 1554 652
rect 1662 648 1666 652
rect 1902 648 1906 652
rect 2366 648 2370 652
rect 2694 648 2698 652
rect 3294 648 3298 652
rect 270 638 274 642
rect 606 638 610 642
rect 694 638 698 642
rect 958 638 962 642
rect 1062 638 1066 642
rect 1198 638 1202 642
rect 1206 638 1210 642
rect 222 628 226 632
rect 398 628 402 632
rect 414 628 418 632
rect 910 628 914 632
rect 1070 628 1074 632
rect 1270 638 1274 642
rect 1422 638 1426 642
rect 1430 638 1434 642
rect 1526 638 1530 642
rect 1558 638 1562 642
rect 1862 638 1866 642
rect 1894 638 1898 642
rect 1926 638 1930 642
rect 1934 638 1938 642
rect 2078 638 2082 642
rect 2126 638 2130 642
rect 2494 638 2498 642
rect 3038 638 3042 642
rect 3198 638 3202 642
rect 3206 638 3210 642
rect 3374 638 3378 642
rect 3390 638 3394 642
rect 1214 628 1218 632
rect 1406 628 1410 632
rect 1462 628 1466 632
rect 1486 628 1490 632
rect 1550 628 1554 632
rect 1678 628 1682 632
rect 1830 628 1834 632
rect 374 618 378 622
rect 430 618 434 622
rect 1094 618 1098 622
rect 1182 618 1186 622
rect 1254 618 1258 622
rect 1358 618 1362 622
rect 1502 618 1506 622
rect 2710 618 2714 622
rect 870 608 874 612
rect 1118 608 1122 612
rect 1270 608 1274 612
rect 1334 608 1338 612
rect 1374 608 1378 612
rect 1942 608 1946 612
rect 2526 608 2530 612
rect 3198 608 3202 612
rect 482 603 486 607
rect 490 603 493 607
rect 493 603 494 607
rect 1514 603 1518 607
rect 1522 603 1525 607
rect 1525 603 1526 607
rect 2538 603 2542 607
rect 2546 603 2549 607
rect 2549 603 2550 607
rect 470 598 474 602
rect 238 588 242 592
rect 574 588 578 592
rect 886 588 890 592
rect 934 588 938 592
rect 1022 588 1026 592
rect 1046 588 1050 592
rect 1054 588 1058 592
rect 3070 588 3074 592
rect 278 578 282 582
rect 686 578 690 582
rect 774 578 778 582
rect 1190 578 1194 582
rect 1958 578 1962 582
rect 1990 578 1994 582
rect 2358 578 2362 582
rect 2422 578 2426 582
rect 2614 578 2618 582
rect 2870 578 2874 582
rect 3102 578 3106 582
rect 182 568 186 572
rect 718 568 722 572
rect 782 568 786 572
rect 910 568 914 572
rect 1310 568 1314 572
rect 1326 568 1330 572
rect 1734 568 1738 572
rect 2638 568 2642 572
rect 302 558 306 562
rect 494 558 498 562
rect 750 558 754 562
rect 934 558 938 562
rect 1006 558 1010 562
rect 1102 558 1106 562
rect 1134 558 1138 562
rect 1166 558 1170 562
rect 1270 558 1274 562
rect 1278 558 1282 562
rect 1422 558 1426 562
rect 1806 558 1810 562
rect 1894 558 1898 562
rect 3094 558 3098 562
rect 110 548 114 552
rect 190 548 194 552
rect 566 548 570 552
rect 606 548 610 552
rect 662 548 666 552
rect 830 548 834 552
rect 854 548 858 552
rect 926 548 930 552
rect 1062 548 1066 552
rect 1110 548 1114 552
rect 1134 548 1138 552
rect 1142 548 1146 552
rect 1158 548 1162 552
rect 1334 548 1338 552
rect 1390 548 1394 552
rect 1406 548 1410 552
rect 598 538 602 542
rect 734 538 738 542
rect 1454 548 1458 552
rect 1486 548 1490 552
rect 1734 548 1738 552
rect 1790 548 1794 552
rect 1918 548 1922 552
rect 1990 548 1994 552
rect 2798 548 2802 552
rect 3166 548 3170 552
rect 3174 548 3178 552
rect 3238 548 3242 552
rect 3294 548 3298 552
rect 886 538 890 542
rect 1078 538 1082 542
rect 1134 538 1138 542
rect 1174 538 1178 542
rect 1190 538 1194 542
rect 1310 538 1314 542
rect 1646 538 1650 542
rect 1718 538 1722 542
rect 1958 538 1962 542
rect 2134 538 2138 542
rect 2670 538 2674 542
rect 2678 538 2682 542
rect 2942 538 2946 542
rect 3014 538 3018 542
rect 3230 538 3234 542
rect 206 528 210 532
rect 222 528 226 532
rect 398 528 402 532
rect 406 528 410 532
rect 798 528 802 532
rect 926 528 930 532
rect 974 528 978 532
rect 1046 528 1050 532
rect 1062 528 1066 532
rect 1542 528 1546 532
rect 1926 528 1930 532
rect 2574 528 2578 532
rect 2814 528 2818 532
rect 3142 528 3146 532
rect 110 518 114 522
rect 278 518 282 522
rect 622 518 626 522
rect 654 518 658 522
rect 766 518 770 522
rect 934 518 938 522
rect 1870 518 1874 522
rect 1950 518 1954 522
rect 2518 518 2522 522
rect 2662 518 2666 522
rect 2670 518 2674 522
rect 2686 518 2690 522
rect 350 508 354 512
rect 614 508 618 512
rect 814 508 818 512
rect 926 508 930 512
rect 1182 508 1186 512
rect 1198 508 1202 512
rect 1406 508 1410 512
rect 1742 508 1746 512
rect 1982 508 1986 512
rect 2198 508 2202 512
rect 2702 508 2706 512
rect 2774 508 2778 512
rect 3086 508 3090 512
rect 3526 508 3530 512
rect 994 503 998 507
rect 1002 503 1005 507
rect 1005 503 1006 507
rect 2026 503 2030 507
rect 2034 503 2037 507
rect 2037 503 2038 507
rect 3042 503 3046 507
rect 3050 503 3053 507
rect 3053 503 3054 507
rect 630 498 634 502
rect 982 498 986 502
rect 1102 498 1106 502
rect 1326 498 1330 502
rect 1334 498 1338 502
rect 1798 498 1802 502
rect 2382 498 2386 502
rect 2766 498 2770 502
rect 3102 498 3106 502
rect 3182 498 3186 502
rect 270 488 274 492
rect 1342 488 1346 492
rect 1822 488 1826 492
rect 1854 488 1858 492
rect 2638 488 2642 492
rect 2734 488 2738 492
rect 3198 488 3202 492
rect 446 478 450 482
rect 470 478 474 482
rect 614 478 618 482
rect 678 478 682 482
rect 870 478 874 482
rect 1150 478 1154 482
rect 1350 478 1354 482
rect 1542 478 1546 482
rect 1846 478 1850 482
rect 2166 478 2170 482
rect 2182 478 2186 482
rect 2326 478 2330 482
rect 2342 478 2346 482
rect 2446 478 2450 482
rect 2638 478 2642 482
rect 2798 478 2802 482
rect 3030 478 3034 482
rect 3222 478 3226 482
rect 3414 478 3418 482
rect 510 468 514 472
rect 582 468 586 472
rect 934 468 938 472
rect 982 468 986 472
rect 1390 468 1394 472
rect 1566 468 1570 472
rect 1886 468 1890 472
rect 2014 468 2018 472
rect 2110 468 2114 472
rect 2174 468 2178 472
rect 2302 468 2306 472
rect 2422 468 2426 472
rect 2598 468 2602 472
rect 2814 468 2818 472
rect 3118 468 3122 472
rect 3318 468 3322 472
rect 3326 468 3330 472
rect 3438 468 3442 472
rect 286 458 290 462
rect 374 458 378 462
rect 406 458 410 462
rect 622 458 626 462
rect 902 458 906 462
rect 1478 458 1482 462
rect 1782 458 1786 462
rect 2390 458 2394 462
rect 3030 458 3034 462
rect 3134 458 3138 462
rect 3142 458 3146 462
rect 3342 458 3346 462
rect 94 448 98 452
rect 862 448 866 452
rect 870 448 874 452
rect 878 448 882 452
rect 1006 448 1010 452
rect 1094 448 1098 452
rect 1118 448 1122 452
rect 1414 448 1418 452
rect 1614 448 1618 452
rect 2174 448 2178 452
rect 2302 448 2306 452
rect 2310 448 2314 452
rect 2694 448 2698 452
rect 2742 448 2746 452
rect 2798 448 2802 452
rect 2902 448 2906 452
rect 2990 448 2994 452
rect 3182 448 3186 452
rect 174 438 178 442
rect 206 438 210 442
rect 238 438 242 442
rect 646 438 650 442
rect 710 438 714 442
rect 950 438 954 442
rect 1054 438 1058 442
rect 1086 438 1090 442
rect 2366 438 2370 442
rect 2790 438 2794 442
rect 2814 438 2818 442
rect 3070 438 3074 442
rect 302 428 306 432
rect 686 428 690 432
rect 1406 428 1410 432
rect 2830 428 2834 432
rect 2950 428 2954 432
rect 3182 428 3186 432
rect 574 418 578 422
rect 1070 418 1074 422
rect 1174 418 1178 422
rect 1550 418 1554 422
rect 1822 418 1826 422
rect 2246 418 2250 422
rect 230 408 234 412
rect 390 408 394 412
rect 510 408 514 412
rect 942 408 946 412
rect 1934 408 1938 412
rect 1942 408 1946 412
rect 3406 408 3410 412
rect 482 403 486 407
rect 490 403 493 407
rect 493 403 494 407
rect 1514 403 1518 407
rect 1522 403 1525 407
rect 1525 403 1526 407
rect 2538 403 2542 407
rect 2546 403 2549 407
rect 2549 403 2550 407
rect 462 398 466 402
rect 598 398 602 402
rect 1022 398 1026 402
rect 1134 398 1138 402
rect 1478 398 1482 402
rect 1630 398 1634 402
rect 1878 398 1882 402
rect 2102 398 2106 402
rect 2278 398 2282 402
rect 2478 398 2482 402
rect 2942 398 2946 402
rect 3430 398 3434 402
rect 414 388 418 392
rect 790 388 794 392
rect 1070 388 1074 392
rect 1078 388 1082 392
rect 1206 388 1210 392
rect 1398 388 1402 392
rect 1870 388 1874 392
rect 3158 388 3162 392
rect 3238 388 3242 392
rect 3326 388 3330 392
rect 358 378 362 382
rect 1542 378 1546 382
rect 1686 378 1690 382
rect 1910 378 1914 382
rect 582 368 586 372
rect 638 368 642 372
rect 678 368 682 372
rect 1446 368 1450 372
rect 1510 368 1514 372
rect 1806 368 1810 372
rect 1966 368 1970 372
rect 2694 368 2698 372
rect 2822 368 2826 372
rect 3038 368 3042 372
rect 270 358 274 362
rect 486 358 490 362
rect 582 358 586 362
rect 614 358 618 362
rect 662 358 666 362
rect 926 358 930 362
rect 1046 358 1050 362
rect 1358 358 1362 362
rect 1630 358 1634 362
rect 1838 358 1842 362
rect 1942 358 1946 362
rect 2214 358 2218 362
rect 2702 358 2706 362
rect 3078 358 3082 362
rect 3430 358 3434 362
rect 70 348 74 352
rect 566 348 570 352
rect 582 348 586 352
rect 694 348 698 352
rect 918 348 922 352
rect 966 348 970 352
rect 1022 348 1026 352
rect 1142 348 1146 352
rect 1158 348 1162 352
rect 1182 348 1186 352
rect 1214 348 1218 352
rect 1270 348 1274 352
rect 1510 348 1514 352
rect 1782 348 1786 352
rect 1814 348 1818 352
rect 1830 348 1834 352
rect 1862 348 1866 352
rect 2102 348 2106 352
rect 2438 348 2442 352
rect 2574 348 2578 352
rect 2590 348 2594 352
rect 2878 348 2882 352
rect 3038 348 3042 352
rect 3078 348 3082 352
rect 3134 348 3138 352
rect 3198 348 3202 352
rect 3478 348 3482 352
rect 542 338 546 342
rect 870 338 874 342
rect 910 338 914 342
rect 1006 338 1010 342
rect 1998 338 2002 342
rect 2126 338 2130 342
rect 2462 338 2466 342
rect 2582 338 2586 342
rect 2822 338 2826 342
rect 2934 338 2938 342
rect 2974 338 2978 342
rect 3102 338 3106 342
rect 3118 338 3122 342
rect 3142 338 3146 342
rect 3230 338 3234 342
rect 3406 338 3410 342
rect 710 328 714 332
rect 1462 328 1466 332
rect 1702 328 1706 332
rect 1798 328 1802 332
rect 2046 328 2050 332
rect 2110 328 2114 332
rect 2270 328 2274 332
rect 2358 328 2362 332
rect 3422 328 3426 332
rect 182 318 186 322
rect 222 318 226 322
rect 398 318 402 322
rect 678 318 682 322
rect 742 318 746 322
rect 774 318 778 322
rect 1710 318 1714 322
rect 2422 318 2426 322
rect 2678 318 2682 322
rect 2974 318 2978 322
rect 3038 318 3042 322
rect 3182 318 3186 322
rect 3262 318 3266 322
rect 1030 308 1034 312
rect 1478 308 1482 312
rect 1678 308 1682 312
rect 1830 308 1834 312
rect 1902 308 1906 312
rect 2006 308 2010 312
rect 2574 308 2578 312
rect 2710 308 2714 312
rect 2774 308 2778 312
rect 2974 308 2978 312
rect 994 303 998 307
rect 1002 303 1005 307
rect 1005 303 1006 307
rect 2026 303 2030 307
rect 2034 303 2037 307
rect 2037 303 2038 307
rect 3042 303 3046 307
rect 3050 303 3053 307
rect 3053 303 3054 307
rect 278 298 282 302
rect 558 298 562 302
rect 830 298 834 302
rect 1110 298 1114 302
rect 1326 298 1330 302
rect 1334 298 1338 302
rect 1926 298 1930 302
rect 2014 298 2018 302
rect 2558 298 2562 302
rect 2614 298 2618 302
rect 2710 298 2714 302
rect 590 288 594 292
rect 1110 288 1114 292
rect 1406 288 1410 292
rect 1430 288 1434 292
rect 1838 288 1842 292
rect 1846 288 1850 292
rect 2318 288 2322 292
rect 2510 288 2514 292
rect 3246 288 3250 292
rect 606 278 610 282
rect 862 278 866 282
rect 934 278 938 282
rect 974 278 978 282
rect 1126 278 1130 282
rect 1142 278 1146 282
rect 1182 278 1186 282
rect 1278 278 1282 282
rect 1462 278 1466 282
rect 1606 278 1610 282
rect 1622 278 1626 282
rect 1694 278 1698 282
rect 1702 278 1706 282
rect 2158 278 2162 282
rect 2398 278 2402 282
rect 2558 278 2562 282
rect 2806 278 2810 282
rect 3006 278 3010 282
rect 3334 278 3338 282
rect 254 268 258 272
rect 614 268 618 272
rect 750 268 754 272
rect 806 268 810 272
rect 1494 268 1498 272
rect 1574 268 1578 272
rect 1582 268 1586 272
rect 1990 268 1994 272
rect 2070 268 2074 272
rect 2142 268 2146 272
rect 2190 268 2194 272
rect 2310 268 2314 272
rect 2334 268 2338 272
rect 2382 268 2386 272
rect 2486 268 2490 272
rect 2502 268 2506 272
rect 2614 268 2618 272
rect 3078 268 3082 272
rect 814 258 818 262
rect 1174 258 1178 262
rect 1374 258 1378 262
rect 1542 258 1546 262
rect 1774 258 1778 262
rect 2294 258 2298 262
rect 2390 258 2394 262
rect 2478 258 2482 262
rect 2686 258 2690 262
rect 2814 258 2818 262
rect 3430 258 3434 262
rect 110 248 114 252
rect 606 248 610 252
rect 630 248 634 252
rect 638 248 642 252
rect 662 248 666 252
rect 750 248 754 252
rect 758 248 762 252
rect 1110 248 1114 252
rect 1262 248 1266 252
rect 1310 248 1314 252
rect 1558 248 1562 252
rect 1622 248 1626 252
rect 1758 248 1762 252
rect 1798 248 1802 252
rect 1830 248 1834 252
rect 2086 248 2090 252
rect 2230 248 2234 252
rect 2302 248 2306 252
rect 2486 248 2490 252
rect 2566 248 2570 252
rect 2798 248 2802 252
rect 1238 238 1242 242
rect 1318 238 1322 242
rect 1550 238 1554 242
rect 1638 238 1642 242
rect 1870 238 1874 242
rect 1974 238 1978 242
rect 1134 228 1138 232
rect 1790 228 1794 232
rect 1918 228 1922 232
rect 1990 238 1994 242
rect 2374 238 2378 242
rect 2718 238 2722 242
rect 1966 228 1970 232
rect 1982 228 1986 232
rect 2710 228 2714 232
rect 2902 228 2906 232
rect 318 218 322 222
rect 518 218 522 222
rect 2326 218 2330 222
rect 2526 218 2530 222
rect 2766 218 2770 222
rect 2990 218 2994 222
rect 30 208 34 212
rect 926 208 930 212
rect 1014 208 1018 212
rect 1022 208 1026 212
rect 1182 208 1186 212
rect 1246 208 1250 212
rect 1254 208 1258 212
rect 1934 208 1938 212
rect 2374 208 2378 212
rect 2486 208 2490 212
rect 3190 208 3194 212
rect 3254 208 3258 212
rect 482 203 486 207
rect 490 203 493 207
rect 493 203 494 207
rect 1514 203 1518 207
rect 1522 203 1525 207
rect 1525 203 1526 207
rect 2538 203 2542 207
rect 2546 203 2549 207
rect 2549 203 2550 207
rect 470 198 474 202
rect 502 198 506 202
rect 878 198 882 202
rect 934 198 938 202
rect 1310 198 1314 202
rect 2270 198 2274 202
rect 2982 198 2986 202
rect 542 188 546 192
rect 2462 188 2466 192
rect 3054 188 3058 192
rect 3094 188 3098 192
rect 1118 178 1122 182
rect 1230 178 1234 182
rect 2174 178 2178 182
rect 2374 178 2378 182
rect 3366 178 3370 182
rect 3390 178 3394 182
rect 190 168 194 172
rect 318 168 322 172
rect 430 168 434 172
rect 446 168 450 172
rect 606 168 610 172
rect 822 168 826 172
rect 830 168 834 172
rect 886 168 890 172
rect 934 168 938 172
rect 1142 168 1146 172
rect 1174 168 1178 172
rect 1414 168 1418 172
rect 1422 168 1426 172
rect 2862 168 2866 172
rect 294 158 298 162
rect 694 158 698 162
rect 702 158 706 162
rect 878 158 882 162
rect 918 158 922 162
rect 958 158 962 162
rect 1166 158 1170 162
rect 2046 158 2050 162
rect 2102 158 2106 162
rect 2142 158 2146 162
rect 2182 158 2186 162
rect 2670 158 2674 162
rect 2678 158 2682 162
rect 2846 158 2850 162
rect 2870 158 2874 162
rect 2902 158 2906 162
rect 2926 158 2930 162
rect 2934 158 2938 162
rect 2950 158 2954 162
rect 2966 158 2970 162
rect 3398 158 3402 162
rect 582 148 586 152
rect 1334 148 1338 152
rect 1342 148 1346 152
rect 1350 148 1354 152
rect 1806 148 1810 152
rect 1870 148 1874 152
rect 2350 148 2354 152
rect 2366 148 2370 152
rect 2414 148 2418 152
rect 2790 148 2794 152
rect 2822 148 2826 152
rect 2886 148 2890 152
rect 2894 148 2898 152
rect 3102 148 3106 152
rect 3110 148 3114 152
rect 3182 148 3186 152
rect 118 138 122 142
rect 214 138 218 142
rect 502 138 506 142
rect 518 138 522 142
rect 622 138 626 142
rect 662 138 666 142
rect 718 138 722 142
rect 734 138 738 142
rect 774 138 778 142
rect 806 138 810 142
rect 838 138 842 142
rect 1118 138 1122 142
rect 1166 138 1170 142
rect 1190 138 1194 142
rect 1230 138 1234 142
rect 1270 138 1274 142
rect 1438 138 1442 142
rect 1454 138 1458 142
rect 1798 138 1802 142
rect 1966 138 1970 142
rect 2406 138 2410 142
rect 2750 138 2754 142
rect 2766 138 2770 142
rect 2942 138 2946 142
rect 3022 138 3026 142
rect 3342 138 3346 142
rect 3366 138 3370 142
rect 3518 138 3522 142
rect 702 128 706 132
rect 758 128 762 132
rect 1078 128 1082 132
rect 1582 128 1586 132
rect 1710 128 1714 132
rect 2062 128 2066 132
rect 2126 128 2130 132
rect 2142 128 2146 132
rect 2398 128 2402 132
rect 2478 128 2482 132
rect 2502 128 2506 132
rect 2590 128 2594 132
rect 2814 128 2818 132
rect 2870 128 2874 132
rect 3070 128 3074 132
rect 3310 128 3314 132
rect 3318 128 3322 132
rect 3350 128 3354 132
rect 3358 128 3362 132
rect 382 118 386 122
rect 446 118 450 122
rect 366 108 370 112
rect 766 118 770 122
rect 894 118 898 122
rect 1302 118 1306 122
rect 1318 118 1322 122
rect 1798 118 1802 122
rect 1806 118 1810 122
rect 2174 118 2178 122
rect 2238 118 2242 122
rect 2486 118 2490 122
rect 2886 118 2890 122
rect 3134 118 3138 122
rect 3302 118 3306 122
rect 3310 118 3314 122
rect 3526 118 3530 122
rect 454 108 458 112
rect 630 108 634 112
rect 878 108 882 112
rect 982 108 986 112
rect 1014 108 1018 112
rect 2166 108 2170 112
rect 2246 108 2250 112
rect 2318 108 2322 112
rect 2326 108 2330 112
rect 2358 108 2362 112
rect 2886 108 2890 112
rect 3014 108 3018 112
rect 3454 108 3458 112
rect 994 103 998 107
rect 1002 103 1005 107
rect 1005 103 1006 107
rect 2026 103 2030 107
rect 2034 103 2037 107
rect 2037 103 2038 107
rect 3042 103 3046 107
rect 3050 103 3053 107
rect 3053 103 3054 107
rect 262 98 266 102
rect 638 98 642 102
rect 822 98 826 102
rect 974 98 978 102
rect 1062 98 1066 102
rect 1798 98 1802 102
rect 2118 98 2122 102
rect 2278 98 2282 102
rect 2326 98 2330 102
rect 2406 98 2410 102
rect 2958 98 2962 102
rect 3030 98 3034 102
rect 3094 98 3098 102
rect 3102 98 3106 102
rect 3326 98 3330 102
rect 3342 98 3346 102
rect 246 88 250 92
rect 398 88 402 92
rect 430 88 434 92
rect 558 88 562 92
rect 566 88 570 92
rect 694 88 698 92
rect 734 88 738 92
rect 782 88 786 92
rect 790 88 794 92
rect 1198 88 1202 92
rect 1246 88 1250 92
rect 2582 88 2586 92
rect 2710 88 2714 92
rect 102 78 106 82
rect 510 78 514 82
rect 942 78 946 82
rect 1022 78 1026 82
rect 1182 78 1186 82
rect 1214 78 1218 82
rect 1286 78 1290 82
rect 1358 78 1362 82
rect 1878 78 1882 82
rect 1902 78 1906 82
rect 1926 78 1930 82
rect 1966 78 1970 82
rect 1990 78 1994 82
rect 2006 78 2010 82
rect 2054 78 2058 82
rect 2686 78 2690 82
rect 2750 78 2754 82
rect 2798 78 2802 82
rect 2886 78 2890 82
rect 422 68 426 72
rect 614 68 618 72
rect 838 68 842 72
rect 862 68 866 72
rect 966 68 970 72
rect 1086 68 1090 72
rect 1142 68 1146 72
rect 1206 68 1210 72
rect 1222 68 1226 72
rect 1294 68 1298 72
rect 1310 68 1314 72
rect 1478 68 1482 72
rect 1494 68 1498 72
rect 3038 78 3042 82
rect 3294 78 3298 82
rect 3438 78 3442 82
rect 3462 78 3466 82
rect 2854 68 2858 72
rect 2862 68 2866 72
rect 2926 68 2930 72
rect 2974 68 2978 72
rect 3030 68 3034 72
rect 3310 68 3314 72
rect 3326 68 3330 72
rect 3342 68 3346 72
rect 3478 68 3482 72
rect 70 58 74 62
rect 230 58 234 62
rect 998 58 1002 62
rect 1102 58 1106 62
rect 1222 58 1226 62
rect 1342 58 1346 62
rect 1358 58 1362 62
rect 1366 58 1370 62
rect 1430 58 1434 62
rect 1446 58 1450 62
rect 1502 58 1506 62
rect 1614 58 1618 62
rect 1630 58 1634 62
rect 2006 58 2010 62
rect 2198 58 2202 62
rect 2222 58 2226 62
rect 2230 58 2234 62
rect 2262 58 2266 62
rect 2334 58 2338 62
rect 2358 58 2362 62
rect 2382 58 2386 62
rect 2782 58 2786 62
rect 3550 58 3554 62
rect 350 48 354 52
rect 478 48 482 52
rect 566 48 570 52
rect 606 48 610 52
rect 662 48 666 52
rect 798 48 802 52
rect 854 48 858 52
rect 1222 48 1226 52
rect 1238 48 1242 52
rect 1454 48 1458 52
rect 1478 48 1482 52
rect 1806 48 1810 52
rect 1902 48 1906 52
rect 2462 48 2466 52
rect 2966 48 2970 52
rect 3142 48 3146 52
rect 3398 48 3402 52
rect 230 38 234 42
rect 390 38 394 42
rect 782 38 786 42
rect 878 38 882 42
rect 1038 38 1042 42
rect 1158 38 1162 42
rect 2294 38 2298 42
rect 2590 38 2594 42
rect 2958 38 2962 42
rect 558 28 562 32
rect 694 28 698 32
rect 710 28 714 32
rect 2574 28 2578 32
rect 2974 38 2978 42
rect 3254 38 3258 42
rect 2966 28 2970 32
rect 598 18 602 22
rect 654 18 658 22
rect 1158 18 1162 22
rect 1214 18 1218 22
rect 1486 18 1490 22
rect 2686 18 2690 22
rect 2766 18 2770 22
rect 2990 18 2994 22
rect 726 8 730 12
rect 814 8 818 12
rect 1054 8 1058 12
rect 1262 8 1266 12
rect 1550 8 1554 12
rect 2342 8 2346 12
rect 2374 8 2378 12
rect 2422 8 2426 12
rect 2758 8 2762 12
rect 2846 8 2850 12
rect 3078 8 3082 12
rect 3334 8 3338 12
rect 482 3 486 7
rect 490 3 493 7
rect 493 3 494 7
rect 1514 3 1518 7
rect 1522 3 1525 7
rect 1525 3 1526 7
rect 2538 3 2542 7
rect 2546 3 2549 7
rect 2549 3 2550 7
<< metal4 >>
rect 992 3303 994 3307
rect 998 3303 1001 3307
rect 1006 3303 1008 3307
rect 2024 3303 2026 3307
rect 2030 3303 2033 3307
rect 2038 3303 2040 3307
rect 3040 3303 3042 3307
rect 3046 3303 3049 3307
rect 3054 3303 3056 3307
rect 690 3298 697 3301
rect 1138 3298 1142 3301
rect 1410 3298 1417 3301
rect 480 3203 482 3207
rect 486 3203 489 3207
rect 494 3203 496 3207
rect 166 3062 169 3068
rect 102 2968 110 2971
rect 6 2652 9 2688
rect 6 2552 9 2558
rect 6 2402 9 2538
rect 14 2471 17 2668
rect 22 2632 25 2668
rect 30 2612 33 2858
rect 46 2842 49 2918
rect 102 2822 105 2968
rect 126 2862 129 2938
rect 138 2908 145 2911
rect 14 2468 22 2471
rect 18 2458 25 2461
rect 22 2372 25 2458
rect 6 2362 9 2368
rect 6 2342 9 2348
rect 30 2342 33 2528
rect 6 2232 9 2268
rect 14 2242 17 2248
rect 38 2242 41 2738
rect 142 2622 145 2908
rect 182 2742 185 2748
rect 62 2452 65 2518
rect 22 2052 25 2168
rect 78 2061 81 2268
rect 86 2072 89 2488
rect 102 2272 105 2448
rect 142 2422 145 2588
rect 154 2518 161 2521
rect 158 2432 161 2518
rect 182 2512 185 2518
rect 198 2502 201 2528
rect 186 2328 193 2331
rect 74 2058 81 2061
rect 78 1982 81 2058
rect 30 1652 33 1858
rect 102 1852 105 1918
rect 6 1042 9 1138
rect 14 1051 17 1298
rect 14 1048 22 1051
rect 6 962 9 978
rect 30 711 33 1648
rect 46 1552 49 1728
rect 38 1548 46 1551
rect 38 1362 41 1548
rect 70 1052 73 1098
rect 86 962 89 1078
rect 58 878 65 881
rect 62 832 65 878
rect 30 708 38 711
rect 30 212 33 708
rect 94 452 97 1438
rect 102 1262 105 1718
rect 110 1512 113 1868
rect 118 1562 121 1958
rect 134 1952 137 2178
rect 118 842 121 858
rect 126 672 129 1828
rect 134 1742 137 1758
rect 134 1281 137 1488
rect 142 1452 145 2058
rect 166 1982 169 2148
rect 174 2142 177 2328
rect 174 2132 177 2138
rect 190 2132 193 2328
rect 206 2182 209 3128
rect 230 2922 233 2948
rect 230 2662 233 2918
rect 238 2872 241 2878
rect 262 2782 265 2948
rect 286 2882 289 2888
rect 278 2852 281 2878
rect 294 2852 297 2858
rect 310 2852 313 3148
rect 606 3082 609 3288
rect 614 3252 617 3258
rect 338 3058 342 3061
rect 570 3058 574 3061
rect 334 3048 342 3051
rect 334 3042 337 3048
rect 370 2868 377 2871
rect 374 2862 377 2868
rect 354 2848 358 2851
rect 282 2828 289 2831
rect 286 2722 289 2828
rect 382 2792 385 3038
rect 406 2898 414 2901
rect 394 2878 398 2881
rect 330 2748 334 2751
rect 350 2718 358 2721
rect 334 2652 337 2668
rect 282 2548 286 2551
rect 214 2492 217 2498
rect 158 1752 161 1958
rect 166 1862 169 1978
rect 174 1851 177 2008
rect 170 1848 177 1851
rect 166 1772 169 1848
rect 158 1652 161 1748
rect 170 1738 174 1741
rect 150 1532 153 1558
rect 158 1522 161 1628
rect 158 1452 161 1518
rect 142 1372 145 1448
rect 134 1278 142 1281
rect 134 1022 137 1138
rect 158 702 161 1448
rect 166 1372 169 1668
rect 182 1652 185 2088
rect 190 1712 193 1888
rect 166 1162 169 1278
rect 174 842 177 1518
rect 182 802 185 938
rect 182 712 185 738
rect 126 662 129 668
rect 182 572 185 708
rect 190 552 193 1598
rect 198 1562 201 1898
rect 206 1572 209 1768
rect 214 1482 217 1948
rect 222 1882 225 1908
rect 230 1862 233 2148
rect 238 2102 241 2198
rect 278 2162 281 2548
rect 294 2471 297 2648
rect 350 2622 353 2718
rect 374 2631 377 2698
rect 406 2692 409 2898
rect 422 2692 425 2868
rect 430 2832 433 2928
rect 386 2638 390 2641
rect 374 2628 385 2631
rect 326 2481 329 2558
rect 370 2518 374 2521
rect 322 2478 329 2481
rect 294 2468 302 2471
rect 286 2371 289 2378
rect 286 2368 294 2371
rect 230 1742 233 1788
rect 238 1742 241 1748
rect 222 1552 225 1658
rect 230 1362 233 1738
rect 238 1712 241 1728
rect 254 1662 257 1778
rect 262 1772 265 2078
rect 270 2072 273 2078
rect 286 1952 289 2208
rect 302 2032 305 2038
rect 310 1981 313 2128
rect 318 2082 321 2168
rect 310 1978 318 1981
rect 270 1611 273 1828
rect 286 1752 289 1918
rect 310 1832 313 1908
rect 334 1862 337 2368
rect 342 2282 345 2328
rect 342 2132 345 2268
rect 278 1682 281 1688
rect 270 1608 278 1611
rect 238 1382 241 1608
rect 246 1392 249 1518
rect 202 1248 206 1251
rect 206 1032 209 1188
rect 206 812 209 1028
rect 198 622 201 648
rect 110 522 113 548
rect 206 442 209 528
rect 178 438 185 441
rect 70 62 73 348
rect 182 322 185 438
rect 110 252 113 268
rect 194 168 198 171
rect 214 142 217 1358
rect 242 1248 246 1251
rect 230 1232 233 1248
rect 226 1058 230 1061
rect 230 922 233 1038
rect 254 942 257 1458
rect 222 532 225 628
rect 238 592 241 858
rect 246 702 249 708
rect 238 542 241 588
rect 246 441 249 508
rect 242 438 249 441
rect 222 408 230 411
rect 222 322 225 408
rect 122 138 126 141
rect 246 92 249 438
rect 254 272 257 908
rect 262 712 265 1458
rect 278 1402 281 1608
rect 286 1602 289 1748
rect 294 1672 297 1798
rect 310 1692 313 1718
rect 318 1712 321 1718
rect 310 1602 313 1668
rect 286 1532 289 1538
rect 294 1462 297 1568
rect 310 1362 313 1418
rect 318 1412 321 1688
rect 326 1602 329 1808
rect 350 1752 353 2368
rect 366 2328 374 2331
rect 366 2322 369 2328
rect 358 1992 361 2268
rect 366 2202 369 2228
rect 366 2171 369 2198
rect 366 2168 374 2171
rect 334 1702 337 1728
rect 350 1692 353 1748
rect 326 1452 329 1568
rect 334 1512 337 1578
rect 330 1428 334 1431
rect 310 1252 313 1358
rect 342 1342 345 1638
rect 358 1532 361 1828
rect 382 1822 385 2628
rect 430 2562 433 2758
rect 438 2652 441 3038
rect 480 3003 482 3007
rect 486 3003 489 3007
rect 494 3003 496 3007
rect 450 2898 457 2901
rect 446 2712 449 2718
rect 454 2702 457 2898
rect 510 2862 513 2868
rect 480 2803 482 2807
rect 486 2803 489 2807
rect 494 2803 496 2807
rect 438 2592 441 2598
rect 434 2518 438 2521
rect 446 2472 449 2688
rect 454 2592 457 2678
rect 454 2502 457 2588
rect 470 2582 473 2798
rect 478 2642 481 2728
rect 498 2708 502 2711
rect 514 2658 518 2661
rect 480 2603 482 2607
rect 486 2603 489 2607
rect 494 2603 496 2607
rect 462 2502 465 2548
rect 526 2542 529 2828
rect 534 2732 537 2738
rect 542 2732 545 3028
rect 554 2878 558 2881
rect 566 2772 569 2788
rect 554 2748 561 2751
rect 542 2642 545 2728
rect 534 2532 537 2548
rect 550 2492 553 2738
rect 558 2652 561 2748
rect 566 2682 569 2768
rect 574 2612 577 2678
rect 582 2581 585 2788
rect 590 2652 593 3048
rect 598 2632 601 3038
rect 606 2642 609 3078
rect 614 3062 617 3088
rect 630 2932 633 3278
rect 574 2578 585 2581
rect 466 2478 470 2481
rect 574 2462 577 2578
rect 582 2542 585 2558
rect 606 2492 609 2638
rect 618 2588 622 2591
rect 630 2572 633 2888
rect 614 2552 617 2558
rect 614 2512 617 2518
rect 598 2452 601 2488
rect 418 2428 422 2431
rect 502 2412 505 2428
rect 390 2342 393 2348
rect 406 2338 414 2341
rect 406 2322 409 2338
rect 410 1978 414 1981
rect 422 1902 425 2308
rect 430 2012 433 2268
rect 438 1982 441 2388
rect 454 2292 457 2338
rect 470 2032 473 2408
rect 480 2403 482 2407
rect 486 2403 489 2407
rect 494 2403 496 2407
rect 502 2222 505 2398
rect 510 2242 513 2428
rect 518 2212 521 2378
rect 526 2331 529 2388
rect 582 2372 585 2428
rect 638 2382 641 2858
rect 654 2801 657 2978
rect 670 2952 673 3288
rect 694 3032 697 3298
rect 710 3268 718 3271
rect 710 3112 713 3268
rect 718 3022 721 3048
rect 726 2892 729 3028
rect 734 2952 737 3228
rect 830 3168 838 3171
rect 758 3002 761 3168
rect 734 2882 737 2948
rect 746 2938 750 2941
rect 798 2932 801 3108
rect 830 3032 833 3168
rect 854 3062 857 3148
rect 814 2942 817 2948
rect 834 2928 838 2931
rect 662 2812 665 2878
rect 734 2872 737 2878
rect 766 2871 769 2928
rect 774 2882 777 2928
rect 846 2922 849 2948
rect 762 2868 769 2871
rect 854 2862 857 2988
rect 886 2982 889 3278
rect 902 3122 905 3148
rect 978 3138 982 3141
rect 902 3082 905 3118
rect 910 3108 918 3111
rect 910 3092 913 3108
rect 992 3103 994 3107
rect 998 3103 1001 3107
rect 1006 3103 1008 3107
rect 1014 3102 1017 3118
rect 942 3052 945 3078
rect 918 2932 921 2938
rect 862 2922 865 2928
rect 906 2868 910 2871
rect 654 2798 665 2801
rect 650 2728 657 2731
rect 654 2722 657 2728
rect 662 2702 665 2798
rect 646 2662 649 2668
rect 646 2642 649 2648
rect 686 2482 689 2798
rect 694 2732 697 2738
rect 718 2652 721 2698
rect 742 2682 745 2718
rect 754 2708 758 2711
rect 774 2652 777 2658
rect 770 2558 774 2561
rect 718 2542 721 2558
rect 658 2458 662 2461
rect 546 2348 553 2351
rect 542 2332 545 2338
rect 526 2328 534 2331
rect 550 2322 553 2348
rect 558 2342 561 2348
rect 574 2342 577 2368
rect 574 2322 577 2338
rect 566 2318 574 2321
rect 480 2203 482 2207
rect 486 2203 489 2207
rect 494 2203 496 2207
rect 502 2162 505 2198
rect 526 2092 529 2238
rect 558 2162 561 2298
rect 566 2262 569 2318
rect 582 2252 585 2368
rect 622 2352 625 2358
rect 654 2352 657 2438
rect 670 2422 673 2458
rect 694 2452 697 2478
rect 594 2318 598 2321
rect 606 2282 609 2318
rect 570 2248 577 2251
rect 574 2242 577 2248
rect 582 2172 585 2248
rect 590 2212 593 2248
rect 546 2158 550 2161
rect 582 2152 585 2158
rect 590 2148 598 2151
rect 602 2148 606 2151
rect 526 2082 529 2088
rect 550 2072 553 2118
rect 530 2068 534 2071
rect 480 2003 482 2007
rect 486 2003 489 2007
rect 494 2003 496 2007
rect 462 1962 465 1998
rect 470 1982 473 1988
rect 398 1752 401 1858
rect 366 1532 369 1718
rect 374 1572 377 1708
rect 398 1622 401 1658
rect 382 1598 390 1601
rect 366 1511 369 1528
rect 362 1508 369 1511
rect 350 1482 353 1498
rect 358 1382 361 1498
rect 350 1322 353 1378
rect 374 1332 377 1558
rect 362 1328 366 1331
rect 298 1248 302 1251
rect 278 732 281 928
rect 286 862 289 1158
rect 362 1068 369 1071
rect 366 992 369 1068
rect 286 842 289 848
rect 270 642 273 668
rect 270 492 273 638
rect 278 582 281 728
rect 286 532 289 838
rect 270 101 273 358
rect 278 302 281 518
rect 286 462 289 528
rect 278 272 281 298
rect 294 162 297 958
rect 306 758 310 761
rect 318 742 321 938
rect 346 858 350 861
rect 334 812 337 858
rect 350 812 353 818
rect 310 692 313 698
rect 334 692 337 808
rect 334 662 337 688
rect 302 652 305 658
rect 302 432 305 558
rect 350 512 353 808
rect 374 732 377 1238
rect 382 962 385 1598
rect 398 1522 401 1558
rect 394 1438 398 1441
rect 406 1302 409 1798
rect 430 1782 433 1948
rect 510 1882 513 2028
rect 530 1978 534 1981
rect 518 1852 521 1878
rect 526 1852 529 1938
rect 542 1932 545 1998
rect 558 1872 561 2138
rect 450 1848 454 1851
rect 414 1662 417 1768
rect 422 1652 425 1668
rect 438 1612 441 1818
rect 480 1803 482 1807
rect 486 1803 489 1807
rect 494 1803 496 1807
rect 414 1572 417 1578
rect 418 1478 422 1481
rect 402 1248 406 1251
rect 390 1182 393 1188
rect 390 962 393 1098
rect 398 972 401 1148
rect 358 382 361 718
rect 374 622 377 668
rect 386 658 393 661
rect 390 652 393 658
rect 382 642 385 648
rect 366 458 374 461
rect 366 452 369 458
rect 390 412 393 648
rect 398 632 401 968
rect 406 621 409 1128
rect 414 952 417 1308
rect 422 1281 425 1468
rect 438 1342 441 1488
rect 446 1482 449 1648
rect 454 1492 457 1768
rect 462 1572 465 1748
rect 494 1742 497 1758
rect 490 1648 494 1651
rect 480 1603 482 1607
rect 486 1603 489 1607
rect 494 1603 496 1607
rect 470 1592 473 1598
rect 446 1392 449 1428
rect 446 1352 449 1388
rect 422 1278 430 1281
rect 422 1072 425 1278
rect 454 1252 457 1348
rect 442 1238 446 1241
rect 462 1202 465 1218
rect 462 1132 465 1158
rect 438 1042 441 1048
rect 470 982 473 1558
rect 502 1542 505 1798
rect 518 1742 521 1848
rect 510 1732 513 1738
rect 518 1672 521 1738
rect 480 1403 482 1407
rect 486 1403 489 1407
rect 494 1403 496 1407
rect 480 1203 482 1207
rect 486 1203 489 1207
rect 494 1203 496 1207
rect 502 1042 505 1348
rect 510 1152 513 1648
rect 518 1362 521 1668
rect 526 1571 529 1778
rect 534 1738 542 1741
rect 534 1592 537 1738
rect 542 1612 545 1708
rect 526 1568 534 1571
rect 530 1538 537 1541
rect 534 1522 537 1538
rect 526 1312 529 1338
rect 518 1062 521 1148
rect 480 1003 482 1007
rect 486 1003 489 1007
rect 494 1003 496 1007
rect 506 978 510 981
rect 470 942 473 958
rect 462 892 465 928
rect 446 842 449 858
rect 462 812 465 848
rect 454 772 457 798
rect 414 632 417 718
rect 406 618 417 621
rect 426 618 430 621
rect 398 532 401 548
rect 406 492 409 528
rect 406 462 409 488
rect 414 392 417 618
rect 438 522 441 708
rect 450 658 457 661
rect 454 642 457 658
rect 450 478 454 481
rect 462 402 465 768
rect 470 682 473 938
rect 480 803 482 807
rect 486 803 489 807
rect 494 803 496 807
rect 470 602 473 658
rect 480 603 482 607
rect 486 603 489 607
rect 494 603 496 607
rect 510 592 513 738
rect 518 682 521 838
rect 526 662 529 1178
rect 534 992 537 1438
rect 542 1192 545 1548
rect 550 1542 553 1548
rect 542 792 545 908
rect 542 722 545 738
rect 498 558 502 561
rect 470 482 473 538
rect 518 502 521 648
rect 550 552 553 1538
rect 558 1402 561 1708
rect 566 1552 569 1968
rect 574 1792 577 2138
rect 590 1991 593 2148
rect 630 2112 633 2168
rect 586 1988 593 1991
rect 598 2062 601 2068
rect 586 1858 590 1861
rect 590 1812 593 1838
rect 574 1541 577 1708
rect 582 1662 585 1738
rect 590 1712 593 1718
rect 590 1551 593 1568
rect 586 1548 593 1551
rect 566 1538 577 1541
rect 566 1372 569 1538
rect 578 1528 582 1531
rect 574 1172 577 1528
rect 582 1092 585 1268
rect 558 852 561 868
rect 566 822 569 1068
rect 582 1041 585 1048
rect 578 1038 585 1041
rect 590 1032 593 1358
rect 574 742 577 888
rect 582 752 585 848
rect 590 832 593 838
rect 558 722 561 728
rect 502 468 510 471
rect 480 403 482 407
rect 486 403 489 407
rect 494 403 496 407
rect 478 361 481 378
rect 478 358 486 361
rect 394 318 398 321
rect 318 172 321 218
rect 454 171 457 318
rect 470 202 473 328
rect 480 203 482 207
rect 486 203 489 207
rect 494 203 496 207
rect 502 202 505 468
rect 450 168 457 171
rect 374 118 382 121
rect 374 112 377 118
rect 266 98 273 101
rect 366 102 369 108
rect 430 92 433 168
rect 502 142 505 198
rect 442 118 446 121
rect 450 108 454 111
rect 390 88 398 91
rect 106 78 110 81
rect 230 42 233 58
rect 350 52 353 88
rect 390 42 393 88
rect 510 82 513 408
rect 542 332 545 338
rect 558 302 561 718
rect 566 552 569 618
rect 566 352 569 548
rect 574 422 577 588
rect 582 472 585 728
rect 590 702 593 798
rect 598 682 601 2058
rect 606 2022 609 2038
rect 606 1742 609 1958
rect 614 1942 617 1948
rect 622 1942 625 2068
rect 622 1872 625 1938
rect 630 1882 633 2078
rect 638 1962 641 2238
rect 646 2112 649 2128
rect 654 2002 657 2348
rect 662 2332 665 2338
rect 674 2238 678 2241
rect 678 2171 681 2198
rect 686 2192 689 2398
rect 694 2232 697 2418
rect 726 2361 729 2408
rect 722 2358 729 2361
rect 702 2172 705 2348
rect 710 2282 713 2348
rect 734 2342 737 2358
rect 734 2321 737 2338
rect 734 2318 742 2321
rect 718 2311 721 2318
rect 718 2308 726 2311
rect 722 2278 726 2281
rect 750 2251 753 2458
rect 758 2442 761 2498
rect 758 2352 761 2368
rect 766 2271 769 2378
rect 762 2268 769 2271
rect 746 2248 753 2251
rect 678 2168 686 2171
rect 690 2078 694 2081
rect 718 2041 721 2068
rect 714 2038 721 2041
rect 638 1882 641 1898
rect 618 1868 622 1871
rect 622 1672 625 1858
rect 646 1812 649 1988
rect 654 1832 657 1988
rect 638 1692 641 1798
rect 670 1761 673 1988
rect 678 1932 681 1958
rect 686 1902 689 1988
rect 726 1982 729 2188
rect 694 1832 697 1908
rect 726 1862 729 1978
rect 686 1772 689 1778
rect 662 1758 673 1761
rect 662 1752 665 1758
rect 646 1742 649 1748
rect 654 1732 657 1738
rect 618 1658 622 1661
rect 606 1562 609 1658
rect 622 1532 625 1658
rect 634 1598 638 1601
rect 610 1528 614 1531
rect 630 1462 633 1508
rect 646 1502 649 1708
rect 654 1702 657 1728
rect 662 1582 665 1608
rect 654 1452 657 1478
rect 606 1162 609 1448
rect 614 1272 617 1278
rect 622 1272 625 1278
rect 622 1092 625 1098
rect 606 1042 609 1068
rect 606 992 609 1038
rect 614 942 617 1068
rect 622 1052 625 1058
rect 630 962 633 1278
rect 622 882 625 938
rect 630 922 633 958
rect 638 892 641 1228
rect 646 1222 649 1348
rect 654 1272 657 1448
rect 670 1312 673 1748
rect 678 1672 681 1678
rect 654 1252 657 1258
rect 662 1112 665 1308
rect 678 1162 681 1638
rect 686 1352 689 1748
rect 694 1682 697 1748
rect 702 1722 705 1768
rect 710 1722 713 1758
rect 710 1582 713 1698
rect 718 1562 721 1748
rect 726 1742 729 1758
rect 726 1712 729 1738
rect 726 1632 729 1638
rect 694 1462 697 1478
rect 686 1162 689 1248
rect 670 1132 673 1138
rect 654 1052 657 1098
rect 654 1042 657 1048
rect 650 948 654 951
rect 606 762 609 828
rect 606 722 609 748
rect 590 652 593 658
rect 598 652 601 678
rect 598 542 601 648
rect 606 632 609 638
rect 606 442 609 548
rect 614 512 617 858
rect 622 822 625 858
rect 662 812 665 1078
rect 670 852 673 1028
rect 654 722 657 788
rect 670 711 673 848
rect 662 708 673 711
rect 586 368 590 371
rect 586 358 590 361
rect 582 342 585 348
rect 518 142 521 218
rect 542 152 545 188
rect 558 92 561 158
rect 582 152 585 338
rect 590 292 593 338
rect 566 92 569 98
rect 426 68 430 71
rect 482 48 486 51
rect 558 51 561 58
rect 558 48 566 51
rect 558 32 561 48
rect 598 22 601 398
rect 606 282 609 438
rect 614 402 617 478
rect 622 462 625 518
rect 630 472 633 498
rect 622 422 625 458
rect 614 362 617 398
rect 638 372 641 708
rect 654 522 657 648
rect 662 552 665 708
rect 678 692 681 948
rect 686 872 689 1158
rect 694 1062 697 1358
rect 702 1152 705 1538
rect 726 1262 729 1318
rect 726 1202 729 1208
rect 734 1152 737 2248
rect 750 2222 753 2248
rect 742 1542 745 1898
rect 750 1752 753 2098
rect 758 2052 761 2238
rect 774 2172 777 2518
rect 782 2342 785 2648
rect 798 2432 801 2678
rect 806 2502 809 2788
rect 814 2532 817 2798
rect 886 2772 889 2868
rect 842 2638 846 2641
rect 846 2602 849 2628
rect 838 2562 841 2568
rect 794 2348 801 2351
rect 782 2332 785 2338
rect 774 2132 777 2138
rect 782 2092 785 2318
rect 798 2312 801 2348
rect 806 2262 809 2468
rect 814 2372 817 2508
rect 834 2458 838 2461
rect 846 2412 849 2418
rect 822 2341 825 2408
rect 818 2338 825 2341
rect 750 1662 753 1748
rect 750 1522 753 1528
rect 742 1402 745 1508
rect 742 1332 745 1398
rect 746 1268 750 1271
rect 746 1198 750 1201
rect 714 1148 718 1151
rect 694 962 697 1058
rect 702 921 705 1148
rect 726 1112 729 1118
rect 710 1062 713 1098
rect 722 1038 726 1041
rect 734 992 737 1038
rect 742 1032 745 1128
rect 742 982 745 1028
rect 702 918 710 921
rect 678 671 681 688
rect 678 668 686 671
rect 670 602 673 668
rect 694 642 697 868
rect 718 862 721 878
rect 714 838 718 841
rect 646 518 654 521
rect 646 442 649 518
rect 686 482 689 578
rect 682 478 686 481
rect 658 358 662 361
rect 606 242 609 248
rect 606 52 609 168
rect 614 72 617 268
rect 622 212 625 328
rect 630 252 633 258
rect 662 252 665 328
rect 678 322 681 368
rect 622 142 625 208
rect 622 108 630 111
rect 622 102 625 108
rect 638 102 641 248
rect 662 152 665 248
rect 686 232 689 428
rect 662 142 665 148
rect 670 51 673 108
rect 686 92 689 228
rect 694 222 697 348
rect 694 162 697 188
rect 702 182 705 838
rect 710 732 713 758
rect 718 712 721 758
rect 726 752 729 918
rect 734 782 737 788
rect 742 702 745 898
rect 722 698 726 701
rect 714 688 718 691
rect 726 652 729 678
rect 710 482 713 648
rect 718 572 721 648
rect 734 552 737 668
rect 750 662 753 1148
rect 758 862 761 2048
rect 790 1991 793 2158
rect 798 2072 801 2138
rect 798 2062 801 2068
rect 790 1988 798 1991
rect 766 1932 769 1978
rect 774 1852 777 1988
rect 774 1772 777 1848
rect 766 1662 769 1688
rect 774 1652 777 1738
rect 782 1682 785 1688
rect 778 1628 782 1631
rect 770 1618 774 1621
rect 778 1578 782 1581
rect 766 1452 769 1498
rect 782 1392 785 1558
rect 782 1262 785 1278
rect 766 1122 769 1248
rect 774 942 777 1088
rect 782 1062 785 1078
rect 782 932 785 998
rect 790 962 793 1778
rect 798 1562 801 1688
rect 798 1252 801 1258
rect 798 1072 801 1158
rect 798 1012 801 1021
rect 758 852 761 858
rect 746 558 750 561
rect 734 542 737 548
rect 710 332 713 438
rect 750 321 753 388
rect 746 318 753 321
rect 742 268 750 271
rect 702 132 705 158
rect 718 142 721 178
rect 742 172 745 268
rect 750 252 753 268
rect 758 252 761 848
rect 766 792 769 798
rect 766 712 769 738
rect 774 692 777 918
rect 782 902 785 918
rect 798 901 801 1008
rect 794 898 801 901
rect 794 888 798 891
rect 798 872 801 878
rect 806 862 809 2258
rect 814 2152 817 2198
rect 822 2092 825 2168
rect 830 2042 833 2358
rect 846 2272 849 2408
rect 814 1692 817 1738
rect 814 1552 817 1688
rect 822 1602 825 1668
rect 822 1492 825 1598
rect 814 1262 817 1468
rect 830 1452 833 1798
rect 838 1482 841 2028
rect 846 2012 849 2268
rect 854 2252 857 2758
rect 870 2752 873 2758
rect 878 2742 881 2758
rect 886 2742 889 2768
rect 870 2631 873 2648
rect 866 2628 873 2631
rect 878 2632 881 2738
rect 878 2582 881 2588
rect 894 2582 897 2698
rect 902 2692 905 2868
rect 926 2752 929 2978
rect 994 2938 998 2941
rect 1014 2932 1017 2948
rect 1002 2928 1006 2931
rect 966 2902 969 2928
rect 974 2922 977 2928
rect 992 2903 994 2907
rect 998 2903 1001 2907
rect 1006 2903 1008 2907
rect 934 2872 937 2888
rect 966 2812 969 2898
rect 950 2762 953 2768
rect 950 2752 953 2758
rect 910 2632 913 2658
rect 870 2332 873 2438
rect 878 2392 881 2468
rect 898 2458 905 2461
rect 878 2362 881 2388
rect 866 2318 873 2321
rect 870 2242 873 2318
rect 854 2171 857 2188
rect 854 2168 862 2171
rect 878 2042 881 2358
rect 886 2352 889 2418
rect 902 2372 905 2458
rect 902 2362 905 2368
rect 910 2351 913 2578
rect 918 2542 921 2698
rect 946 2658 950 2661
rect 946 2638 950 2641
rect 926 2592 929 2628
rect 946 2538 950 2541
rect 910 2348 918 2351
rect 886 2272 889 2338
rect 854 1712 857 1718
rect 822 1162 825 1438
rect 846 1352 849 1688
rect 862 1662 865 1668
rect 870 1662 873 1728
rect 854 1372 857 1588
rect 870 1542 873 1658
rect 862 1512 865 1518
rect 870 1392 873 1408
rect 834 1328 838 1331
rect 850 1308 854 1311
rect 854 1282 857 1288
rect 862 1272 865 1318
rect 870 1302 873 1378
rect 870 1272 873 1278
rect 846 1262 849 1268
rect 850 1228 854 1231
rect 866 1218 870 1221
rect 830 1152 833 1178
rect 838 1152 841 1158
rect 822 1112 825 1148
rect 846 1141 849 1168
rect 846 1138 854 1141
rect 838 1132 841 1138
rect 814 1051 817 1098
rect 814 1048 822 1051
rect 786 798 790 801
rect 790 662 793 748
rect 766 492 769 518
rect 774 492 777 578
rect 782 572 785 638
rect 790 592 793 658
rect 798 532 801 578
rect 774 382 777 488
rect 774 322 777 378
rect 774 142 777 168
rect 722 138 726 141
rect 734 132 737 138
rect 702 92 705 128
rect 734 92 737 128
rect 690 88 694 91
rect 758 82 761 128
rect 766 122 769 138
rect 790 92 793 388
rect 782 82 785 88
rect 798 52 801 308
rect 806 272 809 858
rect 814 742 817 808
rect 822 782 825 968
rect 830 962 833 1058
rect 850 1048 854 1051
rect 838 962 841 1048
rect 862 1012 865 1138
rect 870 1102 873 1128
rect 846 942 849 998
rect 870 992 873 1088
rect 862 942 865 968
rect 870 942 873 968
rect 838 852 841 858
rect 814 512 817 558
rect 822 542 825 778
rect 830 742 833 778
rect 838 742 841 758
rect 830 668 838 671
rect 830 662 833 668
rect 834 548 838 551
rect 846 412 849 938
rect 862 902 865 908
rect 854 752 857 888
rect 870 862 873 868
rect 862 842 865 858
rect 878 852 881 2038
rect 886 1612 889 1988
rect 886 1562 889 1568
rect 886 1522 889 1538
rect 886 1482 889 1488
rect 886 1082 889 1478
rect 878 732 881 738
rect 886 732 889 1048
rect 878 712 881 718
rect 886 702 889 708
rect 854 532 857 548
rect 870 482 873 608
rect 886 592 889 648
rect 878 452 881 518
rect 846 312 849 408
rect 822 298 830 301
rect 806 258 814 261
rect 806 252 809 258
rect 822 172 825 298
rect 862 282 865 448
rect 870 342 873 448
rect 886 432 889 538
rect 878 192 881 198
rect 830 162 833 168
rect 838 142 841 168
rect 878 162 881 188
rect 886 172 889 218
rect 666 48 673 51
rect 702 31 705 38
rect 698 28 705 31
rect 710 32 713 48
rect 786 38 790 41
rect 650 18 654 21
rect 726 12 729 28
rect 806 11 809 138
rect 818 98 822 101
rect 838 72 841 78
rect 846 51 849 158
rect 894 122 897 2268
rect 902 2172 905 2278
rect 902 1952 905 2148
rect 910 2052 913 2088
rect 902 872 905 1748
rect 910 1662 913 1778
rect 910 1532 913 1658
rect 910 1382 913 1398
rect 910 1352 913 1378
rect 910 1132 913 1148
rect 910 1072 913 1098
rect 910 1022 913 1028
rect 910 952 913 998
rect 902 462 905 868
rect 910 692 913 938
rect 910 672 913 688
rect 910 632 913 658
rect 910 572 913 578
rect 910 342 913 358
rect 918 352 921 2338
rect 926 2152 929 2468
rect 934 2352 937 2488
rect 926 2072 929 2108
rect 934 2082 937 2088
rect 942 2012 945 2508
rect 958 2352 961 2768
rect 992 2703 994 2707
rect 998 2703 1001 2707
rect 1006 2703 1008 2707
rect 974 2572 977 2628
rect 998 2532 1001 2688
rect 1006 2522 1009 2538
rect 974 2492 977 2508
rect 992 2503 994 2507
rect 998 2503 1001 2507
rect 1006 2503 1008 2507
rect 966 2392 969 2398
rect 958 2282 961 2348
rect 954 2188 958 2191
rect 950 2052 953 2168
rect 966 2052 969 2308
rect 974 2142 977 2448
rect 1006 2352 1009 2488
rect 1014 2442 1017 2498
rect 1022 2402 1025 3288
rect 1054 3242 1057 3288
rect 1078 3222 1081 3248
rect 1034 3118 1041 3121
rect 1038 2912 1041 3118
rect 1046 2782 1049 2948
rect 1054 2892 1057 2988
rect 1062 2942 1065 2948
rect 1078 2892 1081 3218
rect 1102 3122 1105 3188
rect 1114 3118 1118 3121
rect 1102 3002 1105 3118
rect 1122 3078 1126 3081
rect 1134 3042 1137 3138
rect 1070 2888 1078 2891
rect 1042 2728 1046 2731
rect 1038 2562 1041 2698
rect 1054 2652 1057 2658
rect 1022 2392 1025 2398
rect 992 2303 994 2307
rect 998 2303 1001 2307
rect 1006 2303 1008 2307
rect 982 2292 985 2298
rect 1014 2282 1017 2298
rect 990 2162 993 2168
rect 998 2132 1001 2138
rect 942 1942 945 1948
rect 930 1898 934 1901
rect 926 1832 929 1858
rect 930 1728 937 1731
rect 934 1722 937 1728
rect 942 1711 945 1938
rect 934 1708 945 1711
rect 926 1582 929 1708
rect 926 1532 929 1578
rect 926 1282 929 1458
rect 926 1212 929 1238
rect 934 1142 937 1708
rect 950 1602 953 1928
rect 958 1852 961 1988
rect 942 1542 945 1558
rect 958 1551 961 1788
rect 966 1702 969 1968
rect 982 1942 985 2128
rect 992 2103 994 2107
rect 998 2103 1001 2107
rect 1006 2103 1008 2107
rect 978 1938 982 1941
rect 992 1903 994 1907
rect 998 1903 1001 1907
rect 1006 1903 1008 1907
rect 998 1872 1001 1878
rect 966 1652 969 1688
rect 974 1662 977 1818
rect 986 1768 990 1771
rect 992 1703 994 1707
rect 998 1703 1001 1707
rect 1006 1703 1008 1707
rect 958 1548 969 1551
rect 942 1422 945 1518
rect 958 1402 961 1538
rect 966 1462 969 1548
rect 974 1482 977 1608
rect 1006 1602 1009 1618
rect 982 1512 985 1538
rect 992 1503 994 1507
rect 998 1503 1001 1507
rect 1006 1503 1008 1507
rect 982 1482 985 1498
rect 982 1402 985 1448
rect 946 1368 950 1371
rect 966 1352 969 1368
rect 942 1332 945 1338
rect 942 1262 945 1268
rect 950 1262 953 1328
rect 966 1322 969 1338
rect 974 1312 977 1328
rect 966 1268 974 1271
rect 966 1262 969 1268
rect 982 1262 985 1348
rect 990 1322 993 1448
rect 998 1422 1001 1458
rect 1006 1442 1009 1448
rect 1006 1412 1009 1428
rect 998 1402 1001 1408
rect 1006 1322 1009 1338
rect 992 1303 994 1307
rect 998 1303 1001 1307
rect 1006 1303 1008 1307
rect 942 1192 945 1208
rect 990 1202 993 1208
rect 946 1168 950 1171
rect 958 1161 961 1198
rect 970 1188 974 1191
rect 958 1158 969 1161
rect 926 1132 929 1138
rect 926 852 929 918
rect 934 642 937 1028
rect 942 932 945 1088
rect 950 1062 953 1128
rect 958 982 961 1098
rect 966 1092 969 1158
rect 998 1152 1001 1248
rect 982 1112 985 1118
rect 992 1103 994 1107
rect 998 1103 1001 1107
rect 1006 1103 1008 1107
rect 966 872 969 1068
rect 974 1051 977 1068
rect 990 1052 993 1088
rect 974 1048 982 1051
rect 974 1022 977 1028
rect 974 942 977 998
rect 998 992 1001 1088
rect 1006 1022 1009 1058
rect 982 942 985 958
rect 1006 952 1009 988
rect 982 912 985 918
rect 992 903 994 907
rect 998 903 1001 907
rect 1006 903 1008 907
rect 942 731 945 868
rect 954 858 958 861
rect 982 852 985 898
rect 990 872 993 888
rect 998 872 1001 878
rect 966 782 969 848
rect 974 812 977 838
rect 990 792 993 808
rect 994 758 998 761
rect 942 728 950 731
rect 966 728 974 731
rect 926 552 929 598
rect 934 582 937 588
rect 934 552 937 558
rect 926 512 929 528
rect 934 472 937 518
rect 942 512 945 728
rect 966 691 969 728
rect 958 688 969 691
rect 950 641 953 678
rect 958 662 961 688
rect 950 638 958 641
rect 942 412 945 508
rect 950 442 953 448
rect 958 362 961 638
rect 966 562 969 678
rect 974 642 977 708
rect 992 703 994 707
rect 998 703 1001 707
rect 1006 703 1008 707
rect 982 682 985 698
rect 974 532 977 638
rect 1006 562 1009 578
rect 992 503 994 507
rect 998 503 1001 507
rect 1006 503 1008 507
rect 982 472 985 498
rect 1006 442 1009 448
rect 930 358 934 361
rect 930 278 934 281
rect 926 212 929 228
rect 934 202 937 208
rect 930 168 934 171
rect 950 161 953 178
rect 922 158 929 161
rect 950 158 958 161
rect 866 68 870 71
rect 846 48 854 51
rect 878 42 881 108
rect 926 82 929 158
rect 942 82 945 118
rect 966 72 969 348
rect 1006 342 1009 438
rect 992 303 994 307
rect 998 303 1001 307
rect 1006 303 1008 307
rect 974 102 977 278
rect 1014 212 1017 2148
rect 1022 2032 1025 2358
rect 1030 2342 1033 2538
rect 1054 2532 1057 2608
rect 1062 2522 1065 2878
rect 1070 2852 1073 2888
rect 1038 2472 1041 2498
rect 1038 2362 1041 2448
rect 1038 2282 1041 2358
rect 1022 1752 1025 2018
rect 1022 1522 1025 1708
rect 1030 1672 1033 2038
rect 1038 2022 1041 2278
rect 1046 2092 1049 2348
rect 1054 2061 1057 2398
rect 1062 2352 1065 2488
rect 1070 2462 1073 2828
rect 1086 2752 1089 2898
rect 1086 2562 1089 2568
rect 1078 2542 1081 2558
rect 1062 2272 1065 2278
rect 1070 2202 1073 2368
rect 1062 2062 1065 2078
rect 1054 2058 1062 2061
rect 1046 1922 1049 1968
rect 1038 1712 1041 1728
rect 1046 1721 1049 1758
rect 1054 1732 1057 1908
rect 1078 1832 1081 2488
rect 1086 2342 1089 2508
rect 1094 2452 1097 2948
rect 1118 2901 1121 2968
rect 1114 2898 1121 2901
rect 1126 2912 1129 2938
rect 1118 2882 1121 2888
rect 1126 2862 1129 2908
rect 1142 2892 1145 3148
rect 1150 3012 1153 3078
rect 1150 2992 1153 3008
rect 1182 2932 1185 2948
rect 1110 2762 1113 2788
rect 1102 2728 1110 2731
rect 1102 2492 1105 2728
rect 1110 2561 1113 2688
rect 1126 2662 1129 2668
rect 1134 2572 1137 2868
rect 1198 2752 1201 3158
rect 1186 2748 1190 2751
rect 1146 2668 1153 2671
rect 1150 2632 1153 2668
rect 1158 2662 1161 2668
rect 1174 2602 1177 2728
rect 1214 2682 1217 3078
rect 1230 3022 1233 3288
rect 1246 2992 1249 3248
rect 1286 3242 1289 3258
rect 1230 2942 1233 2968
rect 1262 2892 1265 2908
rect 1286 2882 1289 3158
rect 1294 3082 1297 3298
rect 1338 3138 1342 3141
rect 1318 2922 1321 3038
rect 1298 2888 1302 2891
rect 1326 2852 1329 2928
rect 1238 2752 1241 2848
rect 1226 2748 1230 2751
rect 1226 2698 1230 2701
rect 1110 2558 1118 2561
rect 1130 2548 1137 2551
rect 1118 2512 1121 2548
rect 1134 2532 1137 2548
rect 1150 2541 1153 2568
rect 1146 2538 1153 2541
rect 1126 2528 1134 2531
rect 1102 2472 1105 2478
rect 1114 2448 1121 2451
rect 1118 2442 1121 2448
rect 1118 2292 1121 2298
rect 1086 2082 1089 2198
rect 1094 2062 1097 2258
rect 1106 2218 1110 2221
rect 1102 2072 1105 2118
rect 1086 1932 1089 2028
rect 1094 1872 1097 1878
rect 1062 1772 1065 1778
rect 1046 1718 1057 1721
rect 1038 1672 1041 1688
rect 1046 1552 1049 1708
rect 1054 1672 1057 1718
rect 1062 1672 1065 1678
rect 1054 1662 1057 1668
rect 1054 1582 1057 1588
rect 1054 1552 1057 1558
rect 1030 1512 1033 1538
rect 1026 1468 1030 1471
rect 1054 1462 1057 1538
rect 1062 1482 1065 1508
rect 1022 1442 1025 1458
rect 1030 1452 1033 1458
rect 1062 1442 1065 1448
rect 1022 1382 1025 1398
rect 1030 1351 1033 1408
rect 1026 1348 1033 1351
rect 1022 1342 1025 1348
rect 1030 1332 1033 1338
rect 1038 1321 1041 1378
rect 1046 1352 1049 1418
rect 1030 1318 1041 1321
rect 1030 1301 1033 1318
rect 1022 1298 1033 1301
rect 1022 1252 1025 1298
rect 1030 1272 1033 1288
rect 1022 1202 1025 1208
rect 1022 1152 1025 1158
rect 1030 1112 1033 1258
rect 1038 1252 1041 1308
rect 1038 1212 1041 1228
rect 1046 1182 1049 1328
rect 1054 1232 1057 1418
rect 1062 1262 1065 1378
rect 1070 1322 1073 1768
rect 1078 1392 1081 1798
rect 1086 1742 1089 1788
rect 1094 1782 1097 1808
rect 1086 1452 1089 1558
rect 1094 1422 1097 1708
rect 1102 1582 1105 2018
rect 1118 1972 1121 2278
rect 1126 2242 1129 2528
rect 1134 2442 1137 2448
rect 1134 2372 1137 2438
rect 1146 2378 1153 2381
rect 1162 2378 1166 2381
rect 1150 2372 1153 2378
rect 1134 2282 1137 2328
rect 1142 2262 1145 2338
rect 1150 2292 1153 2308
rect 1126 2142 1129 2218
rect 1142 2152 1145 2258
rect 1166 2252 1169 2338
rect 1174 2262 1177 2548
rect 1182 2281 1185 2428
rect 1190 2332 1193 2438
rect 1182 2278 1190 2281
rect 1158 2142 1161 2248
rect 1178 2228 1182 2231
rect 1198 2092 1201 2408
rect 1206 2312 1209 2658
rect 1214 2552 1217 2558
rect 1222 2512 1225 2518
rect 1214 2342 1217 2448
rect 1230 2412 1233 2668
rect 1246 2502 1249 2818
rect 1254 2572 1257 2758
rect 1318 2712 1321 2808
rect 1326 2712 1329 2718
rect 1302 2602 1305 2638
rect 1254 2492 1257 2548
rect 1278 2532 1281 2538
rect 1242 2458 1246 2461
rect 1214 2312 1217 2318
rect 1230 2281 1233 2368
rect 1246 2312 1249 2348
rect 1254 2342 1257 2488
rect 1262 2482 1265 2488
rect 1286 2458 1294 2461
rect 1286 2452 1289 2458
rect 1270 2382 1273 2388
rect 1270 2352 1273 2378
rect 1294 2372 1297 2438
rect 1278 2302 1281 2368
rect 1226 2278 1233 2281
rect 1230 2122 1233 2278
rect 1238 2192 1241 2288
rect 1250 2268 1254 2271
rect 1110 1602 1113 1738
rect 1118 1711 1121 1828
rect 1134 1802 1137 1948
rect 1142 1842 1145 1858
rect 1126 1732 1129 1778
rect 1134 1732 1137 1768
rect 1118 1708 1126 1711
rect 1118 1582 1121 1668
rect 1134 1642 1137 1648
rect 1130 1618 1134 1621
rect 1134 1602 1137 1608
rect 1086 1372 1089 1378
rect 1078 1302 1081 1318
rect 1054 1142 1057 1228
rect 1070 1202 1073 1268
rect 1078 1242 1081 1268
rect 1086 1262 1089 1338
rect 1094 1272 1097 1368
rect 1102 1312 1105 1498
rect 1118 1432 1121 1488
rect 1126 1452 1129 1578
rect 1142 1572 1145 1778
rect 1150 1762 1153 1978
rect 1158 1872 1161 1878
rect 1158 1712 1161 1728
rect 1166 1712 1169 1988
rect 1182 1902 1185 1948
rect 1206 1882 1209 2118
rect 1254 2042 1257 2118
rect 1262 2082 1265 2288
rect 1278 2282 1281 2298
rect 1286 2292 1289 2308
rect 1294 2282 1297 2308
rect 1294 2132 1297 2148
rect 1206 1871 1209 1878
rect 1206 1868 1214 1871
rect 1166 1672 1169 1678
rect 1182 1662 1185 1798
rect 1206 1722 1209 1728
rect 1198 1712 1201 1718
rect 1194 1678 1198 1681
rect 1170 1658 1174 1661
rect 1142 1552 1145 1568
rect 1150 1532 1153 1608
rect 1174 1602 1177 1618
rect 1154 1518 1158 1521
rect 1166 1512 1169 1558
rect 1174 1531 1177 1598
rect 1198 1572 1201 1588
rect 1174 1528 1182 1531
rect 1206 1522 1209 1718
rect 1214 1662 1217 1828
rect 1222 1571 1225 1838
rect 1246 1772 1249 1968
rect 1254 1942 1257 1948
rect 1270 1802 1273 1888
rect 1278 1872 1281 2038
rect 1286 1942 1289 2108
rect 1294 1931 1297 1988
rect 1302 1952 1305 2468
rect 1310 2092 1313 2268
rect 1310 2022 1313 2068
rect 1294 1928 1302 1931
rect 1254 1782 1257 1788
rect 1242 1738 1246 1741
rect 1222 1568 1230 1571
rect 1134 1452 1137 1488
rect 1118 1322 1121 1348
rect 1090 1248 1094 1251
rect 1102 1242 1105 1258
rect 1110 1242 1113 1278
rect 1110 1192 1113 1218
rect 1118 1192 1121 1318
rect 1126 1252 1129 1388
rect 1142 1342 1145 1468
rect 1150 1402 1153 1418
rect 1158 1392 1161 1398
rect 1150 1312 1153 1328
rect 1158 1322 1161 1328
rect 1062 1132 1065 1158
rect 1030 1082 1033 1088
rect 1022 1062 1025 1068
rect 1038 1061 1041 1078
rect 1034 1058 1041 1061
rect 1054 1062 1057 1098
rect 1022 882 1025 968
rect 1038 942 1041 1048
rect 1054 972 1057 1048
rect 1062 1012 1065 1088
rect 1070 1062 1073 1148
rect 1086 1142 1089 1148
rect 1074 1058 1081 1061
rect 1046 952 1049 958
rect 1054 952 1057 968
rect 1062 942 1065 998
rect 1042 938 1049 941
rect 1038 902 1041 918
rect 1030 872 1033 898
rect 1046 882 1049 938
rect 1054 842 1057 938
rect 1054 832 1057 838
rect 1070 762 1073 998
rect 1078 951 1081 1058
rect 1086 1002 1089 1068
rect 1094 1032 1097 1168
rect 1110 1112 1113 1138
rect 1118 1122 1121 1168
rect 1126 1132 1129 1238
rect 1110 1062 1113 1088
rect 1126 1082 1129 1118
rect 1134 1112 1137 1128
rect 1142 1122 1145 1298
rect 1142 1072 1145 1108
rect 1150 1092 1153 1148
rect 1158 1092 1161 1158
rect 1078 948 1089 951
rect 1078 912 1081 938
rect 1030 672 1033 728
rect 1022 592 1025 658
rect 1030 602 1033 668
rect 1038 642 1041 698
rect 1070 682 1073 698
rect 1078 682 1081 708
rect 1086 682 1089 948
rect 1094 932 1097 1018
rect 1102 962 1105 1018
rect 1110 962 1113 1058
rect 1126 1052 1129 1058
rect 1118 972 1121 1048
rect 1126 962 1129 968
rect 1134 952 1137 1068
rect 1150 972 1153 1068
rect 1142 912 1145 958
rect 1150 912 1153 948
rect 1114 888 1121 891
rect 1118 882 1121 888
rect 1158 882 1161 1058
rect 1166 922 1169 1478
rect 1182 1471 1185 1488
rect 1182 1468 1193 1471
rect 1174 1392 1177 1468
rect 1190 1462 1193 1468
rect 1182 1381 1185 1458
rect 1174 1378 1185 1381
rect 1198 1422 1201 1488
rect 1222 1481 1225 1548
rect 1230 1542 1233 1568
rect 1214 1478 1225 1481
rect 1238 1482 1241 1708
rect 1254 1652 1257 1758
rect 1266 1748 1273 1751
rect 1254 1612 1257 1638
rect 1262 1602 1265 1608
rect 1254 1531 1257 1578
rect 1262 1552 1265 1588
rect 1250 1528 1257 1531
rect 1262 1522 1265 1528
rect 1270 1502 1273 1748
rect 1278 1732 1281 1808
rect 1278 1662 1281 1688
rect 1286 1591 1289 1888
rect 1294 1742 1297 1818
rect 1310 1772 1313 1998
rect 1318 1872 1321 2438
rect 1326 1952 1329 2678
rect 1334 2512 1337 3058
rect 1334 2342 1337 2498
rect 1334 1961 1337 2098
rect 1342 2002 1345 3088
rect 1350 2922 1353 3148
rect 1374 3112 1377 3298
rect 1358 2932 1361 2978
rect 1374 2872 1377 3108
rect 1350 2412 1353 2808
rect 1366 2732 1369 2768
rect 1374 2762 1377 2868
rect 1382 2862 1385 2918
rect 1358 2702 1361 2708
rect 1398 2702 1401 3128
rect 1414 2842 1417 3298
rect 1726 3298 1734 3301
rect 2258 3298 2265 3301
rect 1534 3272 1537 3278
rect 1422 3252 1425 3258
rect 1406 2792 1409 2818
rect 1422 2732 1425 2738
rect 1358 2502 1361 2518
rect 1366 2412 1369 2428
rect 1350 2348 1358 2351
rect 1350 2322 1353 2348
rect 1374 2192 1377 2488
rect 1390 2472 1393 2578
rect 1382 2102 1385 2468
rect 1398 2462 1401 2588
rect 1406 2512 1409 2538
rect 1406 2462 1409 2478
rect 1390 2438 1398 2441
rect 1390 2422 1393 2438
rect 1390 2082 1393 2398
rect 1334 1958 1342 1961
rect 1362 1958 1366 1961
rect 1382 1928 1390 1931
rect 1374 1852 1377 1868
rect 1326 1802 1329 1838
rect 1342 1832 1345 1848
rect 1334 1802 1337 1828
rect 1350 1821 1353 1848
rect 1342 1818 1353 1821
rect 1310 1752 1313 1758
rect 1294 1682 1297 1688
rect 1294 1652 1297 1658
rect 1294 1602 1297 1608
rect 1278 1588 1289 1591
rect 1278 1502 1281 1588
rect 1294 1582 1297 1588
rect 1286 1562 1289 1578
rect 1286 1502 1289 1518
rect 1214 1461 1217 1478
rect 1210 1458 1217 1461
rect 1230 1442 1233 1448
rect 1174 1312 1177 1378
rect 1182 1152 1185 1348
rect 1190 1192 1193 1288
rect 1198 1232 1201 1418
rect 1206 1342 1209 1418
rect 1230 1372 1233 1378
rect 1218 1368 1222 1371
rect 1206 1272 1209 1328
rect 1206 1242 1209 1258
rect 1174 1102 1177 1118
rect 1174 1022 1177 1038
rect 1182 1022 1185 1118
rect 1190 1092 1193 1098
rect 1174 982 1177 1008
rect 1182 992 1185 998
rect 1182 942 1185 968
rect 1182 901 1185 928
rect 1174 898 1185 901
rect 1174 892 1177 898
rect 1110 852 1113 858
rect 1110 712 1113 828
rect 1058 638 1062 641
rect 1046 582 1049 588
rect 1022 402 1025 508
rect 1046 362 1049 528
rect 1054 442 1057 588
rect 1062 532 1065 548
rect 1022 312 1025 348
rect 1030 312 1033 318
rect 1022 262 1025 308
rect 982 112 985 168
rect 1022 112 1025 208
rect 992 103 994 107
rect 998 103 1001 107
rect 1006 103 1008 107
rect 1002 58 1006 61
rect 1014 22 1017 108
rect 1022 82 1025 108
rect 1038 42 1041 48
rect 1054 12 1057 438
rect 1070 422 1073 628
rect 1086 541 1089 588
rect 1082 538 1089 541
rect 1086 442 1089 538
rect 1094 522 1097 618
rect 1118 612 1121 848
rect 1142 832 1145 858
rect 1150 832 1153 878
rect 1166 822 1169 888
rect 1174 852 1177 868
rect 1158 782 1161 788
rect 1134 742 1137 768
rect 1142 702 1145 758
rect 1158 712 1161 748
rect 1134 682 1137 688
rect 1126 672 1129 678
rect 1102 562 1105 598
rect 1110 582 1113 608
rect 1110 552 1113 578
rect 1134 562 1137 578
rect 1142 562 1145 698
rect 1166 692 1169 788
rect 1182 772 1185 868
rect 1178 708 1185 711
rect 1182 702 1185 708
rect 1094 452 1097 518
rect 1102 502 1105 548
rect 1134 542 1137 548
rect 1142 542 1145 548
rect 1062 388 1070 391
rect 1062 102 1065 388
rect 1078 132 1081 388
rect 1110 302 1113 328
rect 1110 282 1113 288
rect 1102 251 1105 258
rect 1102 248 1110 251
rect 1118 182 1121 448
rect 1134 402 1137 538
rect 1150 482 1153 678
rect 1182 652 1185 698
rect 1190 622 1193 1058
rect 1198 1012 1201 1198
rect 1206 1122 1209 1228
rect 1206 1002 1209 1108
rect 1214 1062 1217 1348
rect 1222 1162 1225 1248
rect 1222 1142 1225 1148
rect 1230 1142 1233 1338
rect 1238 1282 1241 1468
rect 1246 1462 1249 1498
rect 1254 1432 1257 1498
rect 1278 1462 1281 1478
rect 1262 1452 1265 1458
rect 1270 1452 1273 1458
rect 1286 1451 1289 1478
rect 1278 1448 1289 1451
rect 1246 1392 1249 1408
rect 1254 1292 1257 1428
rect 1262 1362 1265 1428
rect 1270 1352 1273 1418
rect 1278 1292 1281 1448
rect 1262 1282 1265 1291
rect 1262 1272 1265 1278
rect 1238 1252 1241 1268
rect 1278 1262 1281 1278
rect 1286 1272 1289 1438
rect 1294 1422 1297 1498
rect 1302 1462 1305 1688
rect 1318 1621 1321 1718
rect 1326 1712 1329 1768
rect 1310 1618 1321 1621
rect 1302 1392 1305 1398
rect 1294 1292 1297 1348
rect 1310 1342 1313 1618
rect 1318 1502 1321 1558
rect 1318 1482 1321 1488
rect 1326 1451 1329 1668
rect 1334 1592 1337 1768
rect 1342 1672 1345 1818
rect 1354 1758 1358 1761
rect 1382 1752 1385 1928
rect 1398 1862 1401 2438
rect 1406 2342 1409 2418
rect 1414 2412 1417 2678
rect 1414 2282 1417 2348
rect 1422 2182 1425 2698
rect 1430 2552 1433 3228
rect 1446 3132 1449 3138
rect 1454 3022 1457 3268
rect 1502 3202 1505 3238
rect 1512 3203 1514 3207
rect 1518 3203 1521 3207
rect 1526 3203 1528 3207
rect 1462 3042 1465 3148
rect 1474 3048 1478 3051
rect 1486 3048 1494 3051
rect 1462 2982 1465 3038
rect 1470 2998 1478 3001
rect 1438 2932 1441 2958
rect 1438 2722 1441 2928
rect 1470 2902 1473 2998
rect 1478 2882 1481 2938
rect 1486 2862 1489 3048
rect 1494 3001 1497 3028
rect 1512 3003 1514 3007
rect 1518 3003 1521 3007
rect 1526 3003 1528 3007
rect 1494 2998 1502 3001
rect 1512 2803 1514 2807
rect 1518 2803 1521 2807
rect 1526 2803 1528 2807
rect 1446 2662 1449 2718
rect 1454 2562 1457 2758
rect 1462 2732 1465 2738
rect 1454 2522 1457 2538
rect 1430 2292 1433 2468
rect 1438 2452 1441 2478
rect 1430 2272 1433 2278
rect 1414 2032 1417 2178
rect 1406 1942 1409 1948
rect 1390 1838 1398 1841
rect 1370 1748 1374 1751
rect 1342 1592 1345 1658
rect 1358 1622 1361 1718
rect 1366 1672 1369 1748
rect 1390 1732 1393 1838
rect 1422 1812 1425 2168
rect 1430 1942 1433 2258
rect 1438 2002 1441 2338
rect 1438 1952 1441 1958
rect 1374 1632 1377 1728
rect 1398 1721 1401 1748
rect 1390 1718 1401 1721
rect 1382 1632 1385 1718
rect 1354 1598 1358 1601
rect 1334 1561 1337 1588
rect 1334 1558 1342 1561
rect 1334 1542 1337 1548
rect 1346 1538 1350 1541
rect 1334 1482 1337 1508
rect 1318 1448 1329 1451
rect 1238 1172 1241 1178
rect 1246 1172 1249 1228
rect 1238 1142 1241 1158
rect 1222 992 1225 1108
rect 1230 1052 1233 1088
rect 1246 1071 1249 1148
rect 1254 1142 1257 1198
rect 1262 1122 1265 1188
rect 1254 1112 1257 1118
rect 1270 1082 1273 1168
rect 1246 1068 1254 1071
rect 1198 942 1201 948
rect 1206 932 1209 988
rect 1214 922 1217 948
rect 1206 892 1209 898
rect 1198 792 1201 878
rect 1214 862 1217 898
rect 1206 852 1209 858
rect 1206 802 1209 818
rect 1198 652 1201 738
rect 1206 692 1209 768
rect 1214 681 1217 818
rect 1222 722 1225 948
rect 1230 882 1233 968
rect 1238 932 1241 1048
rect 1246 992 1249 1008
rect 1254 972 1257 1018
rect 1262 962 1265 1068
rect 1250 938 1254 941
rect 1262 922 1265 948
rect 1262 912 1265 918
rect 1238 892 1241 908
rect 1254 892 1257 908
rect 1270 882 1273 1008
rect 1278 972 1281 1238
rect 1286 1182 1289 1218
rect 1294 1152 1297 1258
rect 1302 1222 1305 1318
rect 1310 1272 1313 1278
rect 1318 1262 1321 1448
rect 1326 1252 1329 1338
rect 1334 1332 1337 1468
rect 1342 1442 1345 1528
rect 1350 1422 1353 1498
rect 1342 1362 1345 1368
rect 1342 1322 1345 1348
rect 1310 1248 1318 1251
rect 1302 1162 1305 1198
rect 1310 1152 1313 1248
rect 1318 1192 1321 1238
rect 1334 1221 1337 1298
rect 1342 1262 1345 1268
rect 1334 1218 1342 1221
rect 1334 1192 1337 1198
rect 1318 1162 1321 1168
rect 1294 1112 1297 1148
rect 1302 1142 1305 1148
rect 1286 1042 1289 1108
rect 1294 1082 1297 1098
rect 1302 1081 1305 1128
rect 1310 1092 1313 1148
rect 1334 1142 1337 1178
rect 1326 1122 1329 1128
rect 1322 1108 1329 1111
rect 1302 1078 1313 1081
rect 1294 941 1297 1038
rect 1310 942 1313 1078
rect 1318 1042 1321 1068
rect 1326 1042 1329 1108
rect 1334 1082 1337 1128
rect 1342 1122 1345 1148
rect 1350 1132 1353 1388
rect 1358 1352 1361 1588
rect 1366 1362 1369 1588
rect 1374 1512 1377 1598
rect 1382 1522 1385 1618
rect 1374 1372 1377 1478
rect 1382 1462 1385 1478
rect 1382 1412 1385 1458
rect 1390 1442 1393 1718
rect 1406 1662 1409 1668
rect 1414 1662 1417 1808
rect 1422 1752 1425 1768
rect 1438 1762 1441 1868
rect 1446 1862 1449 2368
rect 1454 2282 1457 2298
rect 1454 2202 1457 2248
rect 1462 2102 1465 2578
rect 1470 2042 1473 2668
rect 1478 2602 1481 2628
rect 1486 2582 1489 2648
rect 1486 2392 1489 2468
rect 1494 2452 1497 2778
rect 1502 2661 1505 2668
rect 1502 2658 1510 2661
rect 1512 2603 1514 2607
rect 1518 2603 1521 2607
rect 1526 2603 1528 2607
rect 1510 2562 1513 2588
rect 1534 2482 1537 3258
rect 1542 2792 1545 3298
rect 1550 2882 1553 2888
rect 1590 2842 1593 2988
rect 1598 2812 1601 3288
rect 1646 3142 1649 3268
rect 1654 3172 1657 3298
rect 1622 3072 1625 3088
rect 1650 2928 1657 2931
rect 1654 2922 1657 2928
rect 1610 2918 1614 2921
rect 1622 2912 1625 2918
rect 1662 2882 1665 3128
rect 1478 1972 1481 2348
rect 1502 2342 1505 2468
rect 1530 2448 1534 2451
rect 1512 2403 1514 2407
rect 1518 2403 1521 2407
rect 1526 2403 1528 2407
rect 1518 2292 1521 2328
rect 1530 2268 1534 2271
rect 1512 2203 1514 2207
rect 1518 2203 1521 2207
rect 1526 2203 1528 2207
rect 1542 2202 1545 2288
rect 1550 2212 1553 2768
rect 1558 2502 1561 2508
rect 1486 1962 1489 2138
rect 1494 2082 1497 2188
rect 1538 2178 1542 2181
rect 1558 2181 1561 2188
rect 1554 2178 1561 2181
rect 1502 2022 1505 2048
rect 1512 2003 1514 2007
rect 1518 2003 1521 2007
rect 1526 2003 1528 2007
rect 1466 1958 1470 1961
rect 1454 1852 1457 1868
rect 1470 1812 1473 1908
rect 1502 1862 1505 1878
rect 1422 1731 1425 1738
rect 1422 1728 1433 1731
rect 1430 1722 1433 1728
rect 1398 1562 1401 1608
rect 1390 1352 1393 1408
rect 1398 1352 1401 1478
rect 1366 1332 1369 1348
rect 1382 1302 1385 1338
rect 1390 1332 1393 1348
rect 1398 1332 1401 1338
rect 1406 1332 1409 1608
rect 1414 1572 1417 1628
rect 1422 1561 1425 1718
rect 1430 1662 1433 1688
rect 1462 1672 1465 1808
rect 1470 1692 1473 1798
rect 1494 1782 1497 1858
rect 1526 1822 1529 1878
rect 1534 1812 1537 1928
rect 1542 1852 1545 1998
rect 1550 1932 1553 1938
rect 1542 1812 1545 1818
rect 1512 1803 1514 1807
rect 1518 1803 1521 1807
rect 1526 1803 1528 1807
rect 1502 1782 1505 1798
rect 1558 1782 1561 2048
rect 1566 2041 1569 2788
rect 1578 2728 1585 2731
rect 1582 2722 1585 2728
rect 1574 2422 1577 2548
rect 1586 2448 1590 2451
rect 1586 2358 1590 2361
rect 1578 2268 1582 2271
rect 1578 2228 1582 2231
rect 1574 2052 1577 2078
rect 1566 2038 1577 2041
rect 1574 1942 1577 2038
rect 1582 1952 1585 2038
rect 1590 1962 1593 2038
rect 1598 2012 1601 2708
rect 1610 2668 1614 2671
rect 1622 2652 1625 2868
rect 1654 2852 1657 2858
rect 1670 2812 1673 3198
rect 1702 3032 1705 3268
rect 1698 2848 1702 2851
rect 1634 2728 1641 2731
rect 1638 2652 1641 2728
rect 1646 2642 1649 2808
rect 1666 2688 1670 2691
rect 1606 2562 1609 2598
rect 1614 2271 1617 2558
rect 1622 2512 1625 2568
rect 1670 2532 1673 2548
rect 1642 2508 1646 2511
rect 1662 2491 1665 2498
rect 1658 2488 1665 2491
rect 1614 2268 1622 2271
rect 1630 2182 1633 2488
rect 1678 2482 1681 2618
rect 1694 2562 1697 2568
rect 1646 2392 1649 2418
rect 1662 2352 1665 2358
rect 1650 2348 1654 2351
rect 1686 2282 1689 2528
rect 1694 2272 1697 2398
rect 1710 2332 1713 3168
rect 1718 2402 1721 3298
rect 1726 3072 1729 3298
rect 1842 3258 1849 3261
rect 1846 3242 1849 3258
rect 1878 3192 1881 3208
rect 1734 2922 1737 2958
rect 1730 2868 1737 2871
rect 1726 2782 1729 2798
rect 1734 2782 1737 2868
rect 1734 2752 1737 2778
rect 1742 2762 1745 3168
rect 1814 3112 1817 3138
rect 1862 3092 1865 3148
rect 1726 2722 1729 2728
rect 1734 2632 1737 2678
rect 1726 2552 1729 2608
rect 1734 2502 1737 2548
rect 1726 2332 1729 2338
rect 1710 2252 1713 2328
rect 1718 2278 1726 2281
rect 1718 2272 1721 2278
rect 1606 2002 1609 2028
rect 1614 1992 1617 2078
rect 1630 2052 1633 2148
rect 1638 2141 1641 2238
rect 1702 2222 1705 2248
rect 1654 2202 1657 2218
rect 1638 2138 1646 2141
rect 1646 2102 1649 2118
rect 1658 2018 1662 2021
rect 1666 1998 1670 2001
rect 1490 1758 1494 1761
rect 1542 1752 1545 1758
rect 1454 1662 1457 1668
rect 1438 1652 1441 1658
rect 1430 1592 1433 1648
rect 1478 1612 1481 1748
rect 1422 1558 1430 1561
rect 1418 1538 1422 1541
rect 1414 1492 1417 1508
rect 1422 1502 1425 1528
rect 1430 1502 1433 1518
rect 1446 1502 1449 1568
rect 1454 1552 1457 1598
rect 1470 1552 1473 1598
rect 1478 1592 1481 1608
rect 1486 1562 1489 1718
rect 1502 1712 1505 1748
rect 1518 1702 1521 1718
rect 1514 1668 1518 1671
rect 1502 1582 1505 1608
rect 1512 1603 1514 1607
rect 1518 1603 1521 1607
rect 1526 1603 1528 1607
rect 1494 1552 1497 1568
rect 1502 1542 1505 1548
rect 1478 1532 1481 1538
rect 1462 1512 1465 1518
rect 1454 1482 1457 1508
rect 1478 1502 1481 1508
rect 1414 1442 1417 1478
rect 1446 1462 1449 1478
rect 1462 1462 1465 1488
rect 1486 1472 1489 1498
rect 1494 1482 1497 1538
rect 1458 1448 1465 1451
rect 1422 1422 1425 1438
rect 1462 1382 1465 1448
rect 1502 1442 1505 1478
rect 1510 1472 1513 1568
rect 1470 1438 1478 1441
rect 1294 938 1302 941
rect 1282 928 1289 931
rect 1230 762 1233 868
rect 1278 832 1281 878
rect 1238 792 1241 828
rect 1286 812 1289 928
rect 1294 928 1302 931
rect 1294 922 1297 928
rect 1294 908 1302 911
rect 1294 852 1297 878
rect 1302 842 1305 898
rect 1310 872 1313 938
rect 1318 902 1321 1018
rect 1334 1012 1337 1068
rect 1326 992 1329 998
rect 1334 922 1337 948
rect 1342 922 1345 1078
rect 1350 1042 1353 1088
rect 1358 992 1361 1268
rect 1366 1252 1369 1288
rect 1366 1072 1369 1138
rect 1374 1082 1377 1258
rect 1390 1232 1393 1318
rect 1382 1142 1385 1168
rect 1390 1142 1393 1178
rect 1318 862 1321 898
rect 1326 868 1334 871
rect 1310 828 1318 831
rect 1246 792 1249 798
rect 1238 751 1241 758
rect 1230 748 1241 751
rect 1230 732 1233 748
rect 1242 728 1246 731
rect 1254 712 1257 798
rect 1262 712 1265 808
rect 1310 802 1313 828
rect 1326 822 1329 868
rect 1342 862 1345 908
rect 1350 832 1353 928
rect 1350 792 1353 828
rect 1286 742 1289 758
rect 1334 742 1337 788
rect 1342 772 1345 778
rect 1350 752 1353 758
rect 1342 742 1345 748
rect 1322 738 1326 741
rect 1358 741 1361 988
rect 1374 932 1377 1068
rect 1398 1052 1401 1288
rect 1414 1232 1417 1318
rect 1422 1262 1425 1298
rect 1430 1262 1433 1268
rect 1422 1242 1425 1248
rect 1406 1102 1409 1158
rect 1422 1131 1425 1218
rect 1430 1192 1433 1208
rect 1438 1172 1441 1348
rect 1470 1332 1473 1438
rect 1510 1432 1513 1468
rect 1518 1462 1521 1568
rect 1526 1532 1529 1578
rect 1534 1562 1537 1598
rect 1542 1522 1545 1658
rect 1550 1612 1553 1728
rect 1566 1702 1569 1928
rect 1574 1792 1577 1798
rect 1582 1762 1585 1948
rect 1622 1922 1625 1938
rect 1630 1922 1633 1928
rect 1590 1851 1593 1868
rect 1598 1862 1601 1898
rect 1626 1858 1630 1861
rect 1590 1848 1598 1851
rect 1578 1738 1582 1741
rect 1590 1732 1593 1818
rect 1574 1691 1577 1728
rect 1598 1722 1601 1838
rect 1606 1822 1609 1838
rect 1606 1732 1609 1788
rect 1614 1721 1617 1798
rect 1606 1718 1617 1721
rect 1566 1688 1577 1691
rect 1550 1552 1553 1598
rect 1558 1571 1561 1668
rect 1566 1582 1569 1688
rect 1558 1568 1569 1571
rect 1534 1442 1537 1458
rect 1542 1452 1545 1458
rect 1550 1452 1553 1528
rect 1558 1482 1561 1518
rect 1566 1471 1569 1568
rect 1574 1562 1577 1578
rect 1582 1572 1585 1648
rect 1590 1572 1593 1668
rect 1606 1662 1609 1718
rect 1614 1658 1622 1661
rect 1614 1632 1617 1658
rect 1590 1552 1593 1558
rect 1598 1552 1601 1618
rect 1606 1562 1609 1618
rect 1630 1592 1633 1828
rect 1638 1792 1641 1858
rect 1646 1732 1649 1928
rect 1654 1852 1657 1878
rect 1662 1872 1665 1958
rect 1670 1952 1673 1958
rect 1670 1922 1673 1948
rect 1670 1802 1673 1868
rect 1678 1791 1681 1958
rect 1694 1881 1697 2058
rect 1702 2012 1705 2038
rect 1710 2002 1713 2068
rect 1718 1962 1721 2178
rect 1726 2062 1729 2068
rect 1734 2062 1737 2448
rect 1750 2402 1753 3068
rect 1782 3052 1785 3058
rect 1818 2938 1822 2941
rect 1766 2922 1769 2938
rect 1794 2928 1798 2931
rect 1758 2702 1761 2718
rect 1758 2582 1761 2698
rect 1742 2342 1745 2348
rect 1746 2328 1750 2331
rect 1758 2302 1761 2578
rect 1766 2562 1769 2918
rect 1786 2848 1790 2851
rect 1774 2812 1777 2848
rect 1774 2652 1777 2808
rect 1794 2768 1798 2771
rect 1790 2712 1793 2738
rect 1774 2562 1777 2568
rect 1782 2542 1785 2558
rect 1790 2492 1793 2608
rect 1734 2032 1737 2038
rect 1726 1972 1729 2028
rect 1742 1942 1745 2158
rect 1754 2098 1758 2101
rect 1766 2082 1769 2488
rect 1782 2362 1785 2378
rect 1774 2342 1777 2348
rect 1782 2332 1785 2358
rect 1790 2202 1793 2208
rect 1774 2072 1777 2168
rect 1782 2138 1790 2141
rect 1766 2042 1769 2058
rect 1690 1878 1697 1881
rect 1694 1861 1697 1868
rect 1718 1862 1721 1928
rect 1742 1872 1745 1928
rect 1734 1862 1737 1868
rect 1690 1858 1697 1861
rect 1706 1858 1710 1861
rect 1750 1852 1753 2028
rect 1782 2022 1785 2138
rect 1798 2132 1801 2588
rect 1806 2202 1809 2798
rect 1814 2141 1817 2898
rect 1830 2832 1833 3068
rect 1862 2932 1865 2988
rect 1862 2922 1865 2928
rect 1878 2912 1881 2928
rect 1846 2882 1849 2888
rect 1842 2858 1846 2861
rect 1866 2768 1870 2771
rect 1830 2622 1833 2688
rect 1838 2602 1841 2618
rect 1846 2592 1849 2748
rect 1878 2612 1881 2908
rect 1890 2878 1894 2881
rect 1902 2862 1905 3048
rect 1910 2912 1913 3148
rect 1918 2862 1921 3298
rect 1926 2902 1929 2928
rect 1918 2702 1921 2858
rect 1926 2802 1929 2808
rect 1862 2582 1865 2598
rect 1822 2491 1825 2558
rect 1834 2538 1841 2541
rect 1838 2532 1841 2538
rect 1846 2522 1849 2528
rect 1822 2488 1830 2491
rect 1834 2328 1838 2331
rect 1830 2308 1838 2311
rect 1830 2292 1833 2308
rect 1846 2152 1849 2198
rect 1814 2138 1822 2141
rect 1846 2141 1849 2148
rect 1842 2138 1849 2141
rect 1790 2122 1793 2128
rect 1774 2012 1777 2018
rect 1774 1952 1777 1978
rect 1758 1882 1761 1938
rect 1782 1932 1785 1948
rect 1802 1928 1806 1931
rect 1766 1902 1769 1918
rect 1774 1892 1777 1928
rect 1794 1908 1798 1911
rect 1710 1848 1718 1851
rect 1670 1788 1681 1791
rect 1654 1722 1657 1788
rect 1654 1682 1657 1688
rect 1638 1582 1641 1608
rect 1558 1468 1569 1471
rect 1558 1441 1561 1468
rect 1542 1438 1561 1441
rect 1494 1362 1497 1408
rect 1502 1402 1505 1418
rect 1512 1403 1514 1407
rect 1518 1403 1521 1407
rect 1526 1403 1528 1407
rect 1534 1352 1537 1408
rect 1542 1321 1545 1438
rect 1566 1421 1569 1458
rect 1534 1318 1545 1321
rect 1550 1418 1569 1421
rect 1414 1128 1425 1131
rect 1430 1132 1433 1168
rect 1406 1032 1409 1048
rect 1414 1012 1417 1128
rect 1422 1032 1425 1118
rect 1438 1062 1441 1098
rect 1446 1082 1449 1238
rect 1454 1182 1457 1188
rect 1462 1172 1465 1268
rect 1470 1232 1473 1268
rect 1478 1262 1481 1288
rect 1462 1152 1465 1158
rect 1470 1122 1473 1168
rect 1478 1152 1481 1208
rect 1486 1132 1489 1288
rect 1494 1192 1497 1208
rect 1512 1203 1514 1207
rect 1518 1203 1521 1207
rect 1526 1203 1528 1207
rect 1486 1092 1489 1098
rect 1350 738 1361 741
rect 1278 728 1286 731
rect 1206 678 1217 681
rect 1206 642 1209 678
rect 1198 632 1201 638
rect 1214 632 1217 638
rect 1178 618 1182 621
rect 1166 562 1169 618
rect 1162 548 1166 551
rect 1174 422 1177 538
rect 1182 512 1185 548
rect 1190 542 1193 578
rect 1158 352 1161 358
rect 1134 348 1142 351
rect 1126 242 1129 278
rect 1134 232 1137 348
rect 1142 262 1145 278
rect 1138 168 1142 171
rect 1166 162 1169 378
rect 1174 348 1182 351
rect 1174 262 1177 348
rect 1182 242 1185 278
rect 1182 212 1185 238
rect 1174 172 1177 178
rect 1110 138 1118 141
rect 1158 138 1166 141
rect 1182 138 1190 141
rect 1090 68 1094 71
rect 1102 62 1105 118
rect 1110 32 1113 138
rect 1142 62 1145 68
rect 1158 42 1161 138
rect 1182 82 1185 138
rect 1198 92 1201 508
rect 1230 412 1233 678
rect 1238 662 1241 698
rect 1278 682 1281 728
rect 1290 708 1297 711
rect 1286 662 1289 668
rect 1294 662 1297 708
rect 1250 658 1257 661
rect 1254 622 1257 658
rect 1270 632 1273 638
rect 1254 432 1257 618
rect 1270 562 1273 608
rect 1278 602 1281 658
rect 1278 542 1281 558
rect 1294 532 1297 558
rect 1302 552 1305 728
rect 1310 612 1313 738
rect 1318 612 1321 688
rect 1330 678 1337 681
rect 1334 672 1337 678
rect 1334 572 1337 608
rect 1322 568 1326 571
rect 1310 562 1313 568
rect 1310 542 1313 548
rect 1206 72 1209 388
rect 1214 352 1217 358
rect 1262 252 1265 428
rect 1270 352 1273 378
rect 1270 278 1278 281
rect 1158 22 1161 38
rect 1214 22 1217 78
rect 1222 72 1225 218
rect 1230 142 1233 178
rect 1226 58 1230 61
rect 1238 52 1241 238
rect 1270 232 1273 278
rect 1246 92 1249 208
rect 1254 192 1257 208
rect 1226 48 1230 51
rect 806 8 814 11
rect 1270 11 1273 138
rect 1286 82 1289 88
rect 1294 72 1297 528
rect 1326 502 1329 538
rect 1334 522 1337 548
rect 1334 502 1337 518
rect 1342 492 1345 678
rect 1350 482 1353 738
rect 1358 622 1361 678
rect 1366 652 1369 918
rect 1390 892 1393 1008
rect 1398 972 1401 1008
rect 1406 962 1409 968
rect 1398 862 1401 958
rect 1422 942 1425 988
rect 1410 928 1414 931
rect 1438 912 1441 988
rect 1422 872 1425 888
rect 1382 858 1390 861
rect 1374 842 1377 848
rect 1382 812 1385 858
rect 1394 848 1398 851
rect 1406 848 1414 851
rect 1406 812 1409 848
rect 1394 808 1401 811
rect 1358 362 1361 618
rect 1374 612 1377 788
rect 1390 702 1393 788
rect 1398 682 1401 808
rect 1430 742 1433 848
rect 1438 842 1441 848
rect 1446 842 1449 1018
rect 1454 982 1457 1078
rect 1462 1072 1465 1078
rect 1462 1032 1465 1038
rect 1470 1002 1473 1038
rect 1478 982 1481 1088
rect 1494 1022 1497 1168
rect 1502 1152 1505 1198
rect 1502 1012 1505 1058
rect 1510 1052 1513 1158
rect 1534 1152 1537 1318
rect 1542 1292 1545 1298
rect 1550 1292 1553 1418
rect 1558 1322 1561 1368
rect 1566 1332 1569 1398
rect 1574 1362 1577 1548
rect 1606 1492 1609 1538
rect 1614 1502 1617 1578
rect 1622 1502 1625 1578
rect 1630 1542 1633 1548
rect 1638 1492 1641 1568
rect 1654 1562 1657 1598
rect 1646 1512 1649 1558
rect 1582 1402 1585 1468
rect 1590 1452 1593 1478
rect 1630 1472 1633 1478
rect 1606 1442 1609 1468
rect 1614 1432 1617 1468
rect 1590 1418 1598 1421
rect 1574 1348 1582 1351
rect 1562 1288 1566 1291
rect 1542 1172 1545 1268
rect 1574 1262 1577 1348
rect 1582 1302 1585 1338
rect 1590 1291 1593 1418
rect 1602 1358 1606 1361
rect 1622 1351 1625 1458
rect 1638 1382 1641 1458
rect 1646 1371 1649 1498
rect 1654 1482 1657 1518
rect 1662 1512 1665 1688
rect 1654 1382 1657 1438
rect 1646 1368 1657 1371
rect 1614 1348 1625 1351
rect 1598 1341 1601 1348
rect 1598 1338 1606 1341
rect 1590 1288 1598 1291
rect 1562 1258 1569 1261
rect 1550 1252 1553 1258
rect 1550 1212 1553 1228
rect 1546 1138 1550 1141
rect 1538 1088 1545 1091
rect 1526 1062 1529 1088
rect 1534 1052 1537 1068
rect 1526 1042 1529 1048
rect 1486 982 1489 1008
rect 1406 732 1409 738
rect 1390 552 1393 578
rect 1390 472 1393 518
rect 1326 292 1329 298
rect 1310 252 1313 268
rect 1314 238 1318 241
rect 1302 102 1305 118
rect 1310 72 1313 198
rect 1334 162 1337 298
rect 1334 152 1337 158
rect 1318 122 1321 138
rect 1342 112 1345 148
rect 1350 92 1353 148
rect 1374 102 1377 258
rect 1390 152 1393 468
rect 1398 392 1401 658
rect 1406 632 1409 638
rect 1406 542 1409 548
rect 1406 512 1409 518
rect 1414 492 1417 738
rect 1454 722 1457 938
rect 1470 892 1473 898
rect 1478 882 1481 978
rect 1494 922 1497 1008
rect 1512 1003 1514 1007
rect 1518 1003 1521 1007
rect 1526 1003 1528 1007
rect 1502 932 1505 998
rect 1478 851 1481 858
rect 1474 848 1481 851
rect 1462 762 1465 848
rect 1478 782 1481 838
rect 1486 762 1489 868
rect 1502 802 1505 868
rect 1510 832 1513 948
rect 1512 803 1514 807
rect 1518 803 1521 807
rect 1526 803 1528 807
rect 1494 732 1497 798
rect 1542 792 1545 1088
rect 1550 972 1553 1098
rect 1558 1082 1561 1228
rect 1566 1202 1569 1258
rect 1582 1172 1585 1288
rect 1590 1212 1593 1288
rect 1558 972 1561 1028
rect 1554 918 1558 921
rect 1558 862 1561 888
rect 1566 862 1569 1148
rect 1574 952 1577 1138
rect 1590 1092 1593 1208
rect 1598 1152 1601 1188
rect 1606 1142 1609 1308
rect 1614 1242 1617 1348
rect 1614 1142 1617 1238
rect 1622 1232 1625 1258
rect 1630 1191 1633 1348
rect 1642 1268 1646 1271
rect 1622 1188 1633 1191
rect 1622 1142 1625 1188
rect 1614 1132 1617 1138
rect 1606 1122 1609 1128
rect 1582 1012 1585 1088
rect 1590 1072 1593 1088
rect 1598 1012 1601 1108
rect 1606 1072 1609 1118
rect 1622 1092 1625 1118
rect 1614 1052 1617 1068
rect 1590 972 1593 1008
rect 1598 962 1601 998
rect 1550 832 1553 848
rect 1574 832 1577 848
rect 1562 828 1569 831
rect 1514 788 1518 791
rect 1438 708 1446 711
rect 1474 708 1478 711
rect 1430 642 1433 678
rect 1438 662 1441 708
rect 1422 632 1425 638
rect 1422 552 1425 558
rect 1422 462 1425 488
rect 1406 292 1409 428
rect 1414 172 1417 448
rect 1438 402 1441 658
rect 1454 652 1457 668
rect 1486 662 1489 718
rect 1466 628 1470 631
rect 1486 622 1489 628
rect 1486 552 1489 598
rect 1454 472 1457 548
rect 1494 482 1497 718
rect 1518 682 1521 698
rect 1506 678 1510 681
rect 1506 668 1510 671
rect 1526 642 1529 688
rect 1542 652 1545 738
rect 1558 712 1561 798
rect 1566 722 1569 828
rect 1574 692 1577 768
rect 1582 732 1585 948
rect 1590 932 1593 958
rect 1614 912 1617 1048
rect 1590 752 1593 858
rect 1606 832 1609 868
rect 1614 772 1617 908
rect 1598 752 1601 758
rect 1622 752 1625 1088
rect 1630 1082 1633 1138
rect 1638 1102 1641 1258
rect 1654 1232 1657 1368
rect 1662 1232 1665 1368
rect 1670 1272 1673 1788
rect 1678 1662 1681 1698
rect 1686 1592 1689 1808
rect 1702 1772 1705 1848
rect 1710 1822 1713 1848
rect 1758 1842 1761 1858
rect 1718 1782 1721 1788
rect 1710 1742 1713 1768
rect 1726 1738 1734 1741
rect 1694 1632 1697 1698
rect 1710 1641 1713 1728
rect 1718 1652 1721 1688
rect 1726 1652 1729 1738
rect 1742 1712 1745 1778
rect 1750 1762 1753 1818
rect 1770 1808 1774 1811
rect 1786 1808 1793 1811
rect 1790 1752 1793 1808
rect 1742 1662 1745 1678
rect 1710 1638 1721 1641
rect 1706 1608 1710 1611
rect 1678 1532 1681 1578
rect 1686 1572 1689 1578
rect 1694 1552 1697 1598
rect 1710 1582 1713 1588
rect 1678 1502 1681 1528
rect 1686 1522 1689 1548
rect 1694 1422 1697 1508
rect 1702 1402 1705 1568
rect 1710 1422 1713 1568
rect 1718 1452 1721 1638
rect 1726 1462 1729 1618
rect 1750 1611 1753 1718
rect 1766 1702 1769 1718
rect 1790 1692 1793 1698
rect 1798 1692 1801 1718
rect 1766 1662 1769 1668
rect 1762 1618 1766 1621
rect 1750 1608 1761 1611
rect 1734 1562 1737 1608
rect 1734 1492 1737 1548
rect 1730 1438 1734 1441
rect 1742 1422 1745 1558
rect 1750 1452 1753 1578
rect 1758 1492 1761 1608
rect 1766 1602 1769 1608
rect 1770 1558 1774 1561
rect 1766 1512 1769 1548
rect 1774 1482 1777 1518
rect 1766 1472 1769 1478
rect 1750 1412 1753 1438
rect 1758 1412 1761 1458
rect 1766 1432 1769 1448
rect 1774 1432 1777 1438
rect 1782 1432 1785 1578
rect 1790 1482 1793 1608
rect 1746 1398 1750 1401
rect 1694 1362 1697 1398
rect 1670 1232 1673 1238
rect 1646 1192 1649 1198
rect 1646 1158 1654 1161
rect 1646 1132 1649 1158
rect 1630 1042 1633 1058
rect 1646 1042 1649 1048
rect 1630 771 1633 968
rect 1638 802 1641 848
rect 1630 768 1638 771
rect 1582 692 1585 698
rect 1550 632 1553 648
rect 1502 612 1505 618
rect 1512 603 1514 607
rect 1518 603 1521 607
rect 1526 603 1528 607
rect 1542 482 1545 528
rect 1458 468 1465 471
rect 1438 371 1441 398
rect 1438 368 1446 371
rect 1462 332 1465 468
rect 1478 402 1481 458
rect 1550 422 1553 608
rect 1512 403 1514 407
rect 1518 403 1521 407
rect 1526 403 1528 407
rect 1510 352 1513 368
rect 1422 172 1425 308
rect 1478 292 1481 308
rect 1430 282 1433 288
rect 1466 278 1470 281
rect 1486 268 1494 271
rect 1438 142 1441 148
rect 1342 78 1358 81
rect 1342 62 1345 78
rect 1354 58 1358 61
rect 1374 61 1377 98
rect 1370 58 1377 61
rect 1430 62 1433 88
rect 1442 58 1446 61
rect 1454 52 1457 138
rect 1478 72 1481 108
rect 1474 48 1478 51
rect 1486 22 1489 268
rect 1542 262 1545 378
rect 1558 252 1561 638
rect 1566 462 1569 468
rect 1590 432 1593 718
rect 1614 682 1617 698
rect 1622 572 1625 718
rect 1646 712 1649 968
rect 1654 742 1657 1138
rect 1662 1122 1665 1128
rect 1670 1112 1673 1158
rect 1666 1068 1670 1071
rect 1666 1048 1673 1051
rect 1670 1022 1673 1048
rect 1662 952 1665 998
rect 1638 538 1646 541
rect 1614 432 1617 448
rect 1630 362 1633 398
rect 1602 278 1606 281
rect 1574 262 1577 268
rect 1512 203 1514 207
rect 1518 203 1521 207
rect 1526 203 1528 207
rect 1494 72 1497 78
rect 1502 62 1505 128
rect 1266 8 1273 11
rect 1550 12 1553 238
rect 1582 132 1585 268
rect 1622 252 1625 278
rect 1638 242 1641 538
rect 1654 442 1657 678
rect 1662 652 1665 948
rect 1670 932 1673 968
rect 1678 962 1681 1338
rect 1686 1332 1689 1348
rect 1694 1332 1697 1338
rect 1718 1322 1721 1398
rect 1758 1342 1761 1398
rect 1766 1342 1769 1348
rect 1726 1328 1734 1331
rect 1754 1328 1758 1331
rect 1686 1201 1689 1258
rect 1694 1212 1697 1318
rect 1702 1302 1705 1318
rect 1714 1298 1718 1301
rect 1702 1232 1705 1268
rect 1710 1232 1713 1258
rect 1686 1198 1697 1201
rect 1686 1132 1689 1148
rect 1694 1092 1697 1198
rect 1702 1122 1705 1158
rect 1710 1102 1713 1188
rect 1718 1172 1721 1288
rect 1726 1202 1729 1328
rect 1734 1262 1737 1308
rect 1750 1302 1753 1308
rect 1758 1272 1761 1288
rect 1742 1192 1745 1258
rect 1766 1242 1769 1328
rect 1774 1302 1777 1418
rect 1782 1302 1785 1308
rect 1778 1278 1782 1281
rect 1790 1281 1793 1398
rect 1798 1392 1801 1578
rect 1806 1552 1809 1848
rect 1814 1722 1817 2128
rect 1846 2102 1849 2118
rect 1854 2102 1857 2518
rect 1870 2372 1873 2588
rect 1878 2372 1881 2378
rect 1886 2371 1889 2638
rect 1894 2542 1897 2568
rect 1902 2562 1905 2668
rect 1886 2368 1894 2371
rect 1910 2322 1913 2618
rect 1918 2612 1921 2618
rect 1862 2112 1865 2318
rect 1894 2292 1897 2308
rect 1822 1962 1825 2078
rect 1886 2072 1889 2198
rect 1910 2182 1913 2258
rect 1894 2122 1897 2178
rect 1902 2062 1905 2178
rect 1918 2132 1921 2528
rect 1858 2048 1862 2051
rect 1834 2028 1838 2031
rect 1830 1982 1833 2008
rect 1838 1922 1841 1998
rect 1846 1922 1849 1988
rect 1854 1952 1857 1958
rect 1830 1902 1833 1918
rect 1854 1852 1857 1938
rect 1862 1922 1865 1968
rect 1878 1962 1881 2058
rect 1902 2051 1905 2058
rect 1898 2048 1905 2051
rect 1910 2052 1913 2078
rect 1918 2012 1921 2088
rect 1926 2072 1929 2138
rect 1926 2002 1929 2028
rect 1934 2022 1937 2928
rect 1942 2852 1945 2858
rect 1950 2762 1953 3218
rect 1958 2852 1961 3198
rect 1990 3122 1993 3128
rect 1966 2822 1969 3108
rect 1986 3048 1990 3051
rect 1966 2672 1969 2738
rect 1982 2702 1985 2898
rect 1998 2871 2001 3298
rect 2162 3288 2166 3291
rect 2178 3288 2185 3291
rect 2182 3272 2185 3288
rect 2034 3258 2038 3261
rect 2024 3103 2026 3107
rect 2030 3103 2033 3107
rect 2038 3103 2040 3107
rect 2010 3088 2014 3091
rect 2062 3062 2065 3148
rect 2170 3128 2174 3131
rect 2158 3078 2166 3081
rect 2050 2948 2054 2951
rect 2026 2938 2030 2941
rect 1994 2868 2001 2871
rect 1994 2858 1998 2861
rect 2002 2728 2006 2731
rect 2006 2691 2009 2708
rect 2014 2702 2017 2928
rect 2024 2903 2026 2907
rect 2030 2903 2033 2907
rect 2038 2903 2040 2907
rect 2078 2892 2081 2928
rect 2086 2922 2089 3078
rect 2098 3068 2102 3071
rect 2062 2732 2065 2758
rect 2070 2742 2073 2748
rect 2024 2703 2026 2707
rect 2030 2703 2033 2707
rect 2038 2703 2040 2707
rect 2002 2688 2009 2691
rect 1998 2608 2006 2611
rect 1982 2422 1985 2538
rect 1942 2332 1945 2338
rect 1950 2332 1953 2358
rect 1874 1928 1881 1931
rect 1890 1928 1897 1931
rect 1830 1772 1833 1848
rect 1822 1722 1825 1738
rect 1830 1682 1833 1748
rect 1838 1742 1841 1798
rect 1846 1752 1849 1768
rect 1854 1762 1857 1848
rect 1870 1842 1873 1848
rect 1862 1831 1865 1838
rect 1862 1828 1873 1831
rect 1870 1812 1873 1828
rect 1878 1772 1881 1928
rect 1886 1872 1889 1908
rect 1894 1892 1897 1928
rect 1918 1922 1921 1928
rect 1926 1882 1929 1958
rect 1846 1672 1849 1728
rect 1838 1668 1846 1671
rect 1806 1402 1809 1528
rect 1822 1522 1825 1668
rect 1814 1452 1817 1478
rect 1822 1382 1825 1488
rect 1830 1452 1833 1558
rect 1838 1512 1841 1668
rect 1846 1552 1849 1658
rect 1826 1368 1830 1371
rect 1798 1292 1801 1298
rect 1790 1278 1801 1281
rect 1778 1228 1782 1231
rect 1742 1162 1745 1188
rect 1750 1182 1753 1188
rect 1718 1122 1721 1148
rect 1734 1142 1737 1158
rect 1718 1098 1726 1101
rect 1702 1092 1705 1098
rect 1710 1072 1713 1098
rect 1718 1082 1721 1098
rect 1686 1022 1689 1038
rect 1694 1012 1697 1048
rect 1686 942 1689 998
rect 1670 862 1673 908
rect 1670 792 1673 848
rect 1670 782 1673 788
rect 1678 632 1681 938
rect 1718 922 1721 1078
rect 1734 1072 1737 1078
rect 1734 952 1737 998
rect 1726 932 1729 948
rect 1750 922 1753 1038
rect 1758 962 1761 1198
rect 1766 1168 1774 1171
rect 1766 1072 1769 1168
rect 1702 912 1705 918
rect 1694 802 1697 878
rect 1702 872 1705 878
rect 1686 782 1689 798
rect 1710 792 1713 918
rect 1742 892 1745 908
rect 1750 892 1753 898
rect 1726 862 1729 878
rect 1758 802 1761 808
rect 1766 782 1769 1048
rect 1774 772 1777 1148
rect 1782 942 1785 1158
rect 1790 1132 1793 1228
rect 1798 1142 1801 1278
rect 1806 1252 1809 1338
rect 1806 1162 1809 1248
rect 1814 1182 1817 1358
rect 1822 1322 1825 1348
rect 1822 1282 1825 1298
rect 1830 1212 1833 1338
rect 1838 1282 1841 1488
rect 1846 1422 1849 1548
rect 1846 1402 1849 1408
rect 1846 1372 1849 1378
rect 1846 1332 1849 1358
rect 1846 1252 1849 1268
rect 1854 1252 1857 1758
rect 1862 1752 1865 1768
rect 1870 1722 1873 1768
rect 1862 1592 1865 1718
rect 1886 1682 1889 1848
rect 1894 1842 1897 1848
rect 1878 1662 1881 1678
rect 1870 1582 1873 1618
rect 1862 1322 1865 1548
rect 1870 1472 1873 1578
rect 1878 1562 1881 1648
rect 1894 1572 1897 1828
rect 1902 1702 1905 1868
rect 1910 1842 1913 1848
rect 1910 1828 1918 1831
rect 1910 1762 1913 1828
rect 1926 1812 1929 1858
rect 1934 1832 1937 1998
rect 1942 1952 1945 2018
rect 1950 2012 1953 2318
rect 1958 2292 1961 2318
rect 1966 2282 1969 2358
rect 1998 2352 2001 2608
rect 2014 2571 2017 2598
rect 2010 2568 2017 2571
rect 2038 2532 2041 2608
rect 2024 2503 2026 2507
rect 2030 2503 2033 2507
rect 2038 2503 2040 2507
rect 2046 2502 2049 2548
rect 2006 2472 2009 2488
rect 2006 2312 2009 2328
rect 2014 2272 2017 2318
rect 2024 2303 2026 2307
rect 2030 2303 2033 2307
rect 2038 2303 2040 2307
rect 2046 2302 2049 2398
rect 2022 2262 2025 2278
rect 2054 2172 2057 2648
rect 2062 2522 2065 2528
rect 2070 2502 2073 2538
rect 2066 2468 2073 2471
rect 2070 2342 2073 2468
rect 2070 2262 2073 2268
rect 2078 2201 2081 2858
rect 2086 2732 2089 2918
rect 2110 2872 2113 2878
rect 2102 2672 2105 2768
rect 2118 2732 2121 2908
rect 2126 2812 2129 3048
rect 2122 2718 2126 2721
rect 2118 2668 2126 2671
rect 2118 2662 2121 2668
rect 2134 2572 2137 2728
rect 2142 2642 2145 2648
rect 2134 2502 2137 2568
rect 2150 2492 2153 2868
rect 2158 2822 2161 3078
rect 2178 3068 2182 3071
rect 2182 2952 2185 3058
rect 2190 3042 2193 3138
rect 2198 2952 2201 3298
rect 2234 3288 2238 3291
rect 2214 3252 2217 3258
rect 2222 3122 2225 3138
rect 2206 3102 2209 3108
rect 2214 3092 2217 3108
rect 2178 2948 2182 2951
rect 2210 2858 2214 2861
rect 2182 2802 2185 2828
rect 2122 2358 2126 2361
rect 2098 2348 2102 2351
rect 2098 2328 2105 2331
rect 2102 2322 2105 2328
rect 2074 2198 2081 2201
rect 2086 2202 2089 2218
rect 2062 2182 2065 2198
rect 2086 2172 2089 2198
rect 2094 2162 2097 2268
rect 2102 2172 2105 2288
rect 2110 2282 2113 2348
rect 2110 2272 2113 2278
rect 2134 2272 2137 2488
rect 2146 2278 2150 2281
rect 2126 2252 2129 2268
rect 1958 2142 1961 2148
rect 2046 2112 2049 2128
rect 2024 2103 2026 2107
rect 2030 2103 2033 2107
rect 2038 2103 2040 2107
rect 2054 2051 2057 2098
rect 2062 2062 2065 2078
rect 2094 2062 2097 2148
rect 2134 2102 2137 2118
rect 2054 2048 2062 2051
rect 1942 1872 1945 1928
rect 1934 1802 1937 1808
rect 1926 1772 1929 1778
rect 1918 1751 1921 1768
rect 1910 1748 1921 1751
rect 1910 1652 1913 1748
rect 1934 1741 1937 1778
rect 1942 1762 1945 1768
rect 1930 1738 1937 1741
rect 1886 1562 1889 1568
rect 1886 1522 1889 1538
rect 1878 1492 1881 1508
rect 1894 1502 1897 1538
rect 1886 1492 1889 1498
rect 1902 1462 1905 1598
rect 1870 1392 1873 1398
rect 1894 1382 1897 1398
rect 1910 1382 1913 1518
rect 1894 1362 1897 1368
rect 1874 1358 1878 1361
rect 1878 1332 1881 1348
rect 1886 1332 1889 1348
rect 1862 1282 1865 1308
rect 1838 1212 1841 1218
rect 1802 1128 1806 1131
rect 1814 1122 1817 1138
rect 1806 1102 1809 1108
rect 1798 962 1801 1098
rect 1806 942 1809 1088
rect 1790 938 1798 941
rect 1722 748 1726 751
rect 1734 742 1737 748
rect 1782 742 1785 848
rect 1790 802 1793 938
rect 1798 902 1801 908
rect 1798 802 1801 888
rect 1814 872 1817 1088
rect 1822 1062 1825 1158
rect 1830 1092 1833 1108
rect 1838 1082 1841 1208
rect 1846 1102 1849 1238
rect 1854 1142 1857 1248
rect 1870 1212 1873 1218
rect 1878 1201 1881 1318
rect 1886 1221 1889 1298
rect 1894 1272 1897 1358
rect 1902 1302 1905 1318
rect 1910 1292 1913 1368
rect 1918 1362 1921 1678
rect 1926 1662 1929 1728
rect 1950 1692 1953 1898
rect 1958 1782 1961 2018
rect 1998 1982 2001 2048
rect 1974 1932 1977 1968
rect 1990 1912 1993 1968
rect 1998 1948 2006 1951
rect 1998 1922 2001 1948
rect 2038 1922 2041 1928
rect 2046 1912 2049 1968
rect 2086 1962 2089 2058
rect 2130 2048 2134 2051
rect 2142 2002 2145 2058
rect 2150 2052 2153 2078
rect 2158 2071 2161 2638
rect 2166 2292 2169 2758
rect 2190 2552 2193 2748
rect 2178 2528 2182 2531
rect 2198 2412 2201 2568
rect 2206 2562 2209 2828
rect 2222 2722 2225 3078
rect 2238 2681 2241 2988
rect 2246 2982 2249 3288
rect 2262 3132 2265 3298
rect 2630 3298 2638 3301
rect 3082 3298 3089 3301
rect 2310 3262 2313 3268
rect 2310 3052 2313 3138
rect 2370 3108 2374 3111
rect 2318 3042 2321 3088
rect 2438 3072 2441 3078
rect 2250 2868 2254 2871
rect 2238 2678 2246 2681
rect 2218 2638 2225 2641
rect 2206 2522 2209 2528
rect 2166 2272 2169 2278
rect 2194 2268 2198 2271
rect 2206 2262 2209 2268
rect 2174 2232 2177 2248
rect 2182 2112 2185 2168
rect 2214 2102 2217 2628
rect 2222 2622 2225 2638
rect 2166 2082 2169 2088
rect 2206 2082 2209 2088
rect 2222 2082 2225 2598
rect 2230 2352 2233 2368
rect 2238 2132 2241 2168
rect 2158 2068 2169 2071
rect 2014 1871 2017 1908
rect 2024 1903 2026 1907
rect 2030 1903 2033 1907
rect 2038 1903 2040 1907
rect 2014 1868 2025 1871
rect 2022 1862 2025 1868
rect 1990 1852 1993 1858
rect 1998 1848 2006 1851
rect 2014 1851 2017 1858
rect 2014 1848 2022 1851
rect 1998 1842 2001 1848
rect 1994 1798 1998 1801
rect 1958 1702 1961 1758
rect 1982 1712 1985 1728
rect 1990 1692 1993 1748
rect 2022 1732 2025 1828
rect 2038 1772 2041 1838
rect 2046 1738 2054 1741
rect 1938 1688 1942 1691
rect 1938 1668 1945 1671
rect 1934 1532 1937 1548
rect 1942 1522 1945 1668
rect 1958 1662 1961 1668
rect 1966 1592 1969 1668
rect 1986 1658 1990 1661
rect 1998 1652 2001 1698
rect 1950 1552 1953 1588
rect 1926 1482 1929 1498
rect 1934 1471 1937 1498
rect 1926 1468 1937 1471
rect 1926 1352 1929 1468
rect 1934 1352 1937 1438
rect 1942 1412 1945 1428
rect 1942 1352 1945 1358
rect 1938 1318 1945 1321
rect 1902 1271 1905 1288
rect 1902 1268 1910 1271
rect 1886 1218 1894 1221
rect 1870 1198 1881 1201
rect 1870 1182 1873 1198
rect 1838 932 1841 958
rect 1846 942 1849 958
rect 1854 942 1857 1138
rect 1862 982 1865 1158
rect 1886 1152 1889 1168
rect 1870 972 1873 1148
rect 1878 1112 1881 1128
rect 1886 1122 1889 1128
rect 1826 928 1830 931
rect 1846 858 1862 861
rect 1846 852 1849 858
rect 1826 848 1830 851
rect 1870 822 1873 948
rect 1878 922 1881 1068
rect 1886 942 1889 1118
rect 1894 1102 1897 1188
rect 1894 1062 1897 1078
rect 1902 1062 1905 1258
rect 1910 1212 1913 1258
rect 1918 1222 1921 1298
rect 1902 1042 1905 1048
rect 1702 652 1705 668
rect 1710 662 1713 688
rect 1726 682 1729 738
rect 1782 702 1785 728
rect 1790 712 1793 798
rect 1830 742 1833 758
rect 1842 748 1846 751
rect 1854 722 1857 738
rect 1734 652 1737 688
rect 1758 662 1761 688
rect 1782 672 1785 678
rect 1766 662 1769 668
rect 1790 662 1793 668
rect 1734 552 1737 568
rect 1718 532 1721 538
rect 1742 482 1745 508
rect 1778 458 1782 461
rect 1678 282 1681 308
rect 1686 281 1689 378
rect 1778 348 1782 351
rect 1702 332 1705 348
rect 1686 278 1694 281
rect 1686 272 1689 278
rect 1702 272 1705 278
rect 1710 132 1713 318
rect 1758 252 1761 268
rect 1770 258 1774 261
rect 1790 232 1793 548
rect 1798 512 1801 698
rect 1826 688 1830 691
rect 1814 682 1817 688
rect 1810 558 1814 561
rect 1798 332 1801 498
rect 1822 492 1825 658
rect 1854 652 1857 658
rect 1862 642 1865 748
rect 1870 692 1873 698
rect 1830 502 1833 628
rect 1878 622 1881 918
rect 1894 912 1897 1008
rect 1910 992 1913 1058
rect 1918 982 1921 1178
rect 1926 1172 1929 1318
rect 1942 1312 1945 1318
rect 1942 1271 1945 1288
rect 1938 1268 1945 1271
rect 1950 1262 1953 1328
rect 1942 1192 1945 1258
rect 1934 1132 1937 1148
rect 1926 1062 1929 1108
rect 1934 1082 1937 1108
rect 1942 1052 1945 1128
rect 1950 1072 1953 1178
rect 1958 1132 1961 1578
rect 2006 1572 2009 1678
rect 2014 1582 2017 1708
rect 2024 1703 2026 1707
rect 2030 1703 2033 1707
rect 2038 1703 2040 1707
rect 2046 1652 2049 1738
rect 2062 1732 2065 1958
rect 2094 1951 2097 1968
rect 2094 1948 2102 1951
rect 2070 1832 2073 1838
rect 2070 1802 2073 1828
rect 2054 1642 2057 1708
rect 2078 1682 2081 1848
rect 2086 1792 2089 1808
rect 2094 1782 2097 1938
rect 2110 1932 2113 1998
rect 2110 1762 2113 1858
rect 2118 1772 2121 1858
rect 2086 1692 2089 1748
rect 2126 1732 2129 1918
rect 2166 1912 2169 2068
rect 2186 2058 2190 2061
rect 2246 2051 2249 2668
rect 2258 2528 2262 2531
rect 2270 2521 2273 3018
rect 2286 2752 2289 2858
rect 2350 2712 2353 3058
rect 2366 2932 2369 2948
rect 2342 2682 2345 2698
rect 2310 2672 2313 2678
rect 2350 2552 2353 2698
rect 2262 2518 2273 2521
rect 2254 2462 2257 2478
rect 2254 2162 2257 2178
rect 2262 2052 2265 2518
rect 2270 2332 2273 2338
rect 2246 2048 2257 2051
rect 2198 1982 2201 2038
rect 2154 1908 2158 1911
rect 2158 1862 2161 1898
rect 2134 1742 2137 1748
rect 2118 1712 2121 1718
rect 2134 1692 2137 1728
rect 2054 1572 2057 1588
rect 1966 1402 1969 1568
rect 2062 1562 2065 1598
rect 2010 1558 2017 1561
rect 2042 1558 2046 1561
rect 1966 1342 1969 1378
rect 1974 1331 1977 1548
rect 1982 1532 1985 1538
rect 1990 1492 1993 1558
rect 2006 1512 2009 1518
rect 2014 1512 2017 1558
rect 2070 1552 2073 1678
rect 2102 1652 2105 1678
rect 2110 1672 2113 1678
rect 2118 1648 2126 1651
rect 2024 1503 2026 1507
rect 2030 1503 2033 1507
rect 2038 1503 2040 1507
rect 2046 1502 2049 1548
rect 2054 1542 2057 1548
rect 2094 1542 2097 1588
rect 2110 1582 2113 1638
rect 2118 1622 2121 1648
rect 2006 1482 2009 1498
rect 1990 1372 1993 1478
rect 2030 1432 2033 1448
rect 1966 1328 1977 1331
rect 1966 1172 1969 1328
rect 1982 1322 1985 1348
rect 1974 1292 1977 1298
rect 1982 1222 1985 1268
rect 1990 1242 1993 1338
rect 1958 1042 1961 1108
rect 1966 1042 1969 1108
rect 1974 1071 1977 1218
rect 1998 1182 2001 1428
rect 2006 1332 2009 1408
rect 2030 1372 2033 1418
rect 2014 1302 2017 1358
rect 2030 1322 2033 1348
rect 2038 1342 2041 1468
rect 2046 1391 2049 1498
rect 2054 1432 2057 1538
rect 2102 1532 2105 1538
rect 2118 1532 2121 1558
rect 2054 1402 2057 1408
rect 2046 1388 2057 1391
rect 2046 1332 2049 1358
rect 2054 1352 2057 1388
rect 2046 1312 2049 1318
rect 2054 1312 2057 1348
rect 2024 1303 2026 1307
rect 2030 1303 2033 1307
rect 2038 1303 2040 1307
rect 2014 1282 2017 1298
rect 1982 1152 1985 1158
rect 1986 1138 1993 1141
rect 1990 1122 1993 1138
rect 1974 1068 1982 1071
rect 1902 952 1905 978
rect 1886 908 1894 911
rect 1886 672 1889 908
rect 1910 822 1913 838
rect 1918 832 1921 908
rect 1926 872 1929 948
rect 1934 912 1937 1038
rect 1990 1022 1993 1108
rect 1950 942 1953 968
rect 1958 952 1961 968
rect 1970 948 1974 951
rect 1942 921 1945 938
rect 1942 918 1950 921
rect 1970 918 1974 921
rect 1950 891 1953 898
rect 1982 892 1985 988
rect 1998 982 2001 1148
rect 2006 1102 2009 1168
rect 1950 888 1958 891
rect 1942 882 1945 888
rect 1930 848 1934 851
rect 1846 482 1849 618
rect 1874 518 1881 521
rect 1806 292 1809 368
rect 1822 351 1825 418
rect 1838 352 1841 358
rect 1822 348 1830 351
rect 1814 282 1817 348
rect 1830 292 1833 308
rect 1838 292 1841 308
rect 1854 291 1857 488
rect 1878 402 1881 518
rect 1886 472 1889 658
rect 1894 642 1897 818
rect 1902 782 1905 788
rect 1934 722 1937 748
rect 1894 562 1897 598
rect 1866 388 1870 391
rect 1850 288 1857 291
rect 1862 282 1865 348
rect 1902 312 1905 648
rect 1910 382 1913 678
rect 1926 642 1929 658
rect 1934 642 1937 648
rect 1918 552 1921 618
rect 1942 612 1945 858
rect 1966 851 1969 868
rect 1962 848 1969 851
rect 1990 762 1993 828
rect 1962 738 1966 741
rect 1950 732 1953 738
rect 1918 432 1921 438
rect 1806 251 1809 268
rect 1802 248 1809 251
rect 1822 248 1830 251
rect 1822 242 1825 248
rect 1870 152 1873 238
rect 1918 232 1921 428
rect 1926 302 1929 528
rect 1950 522 1953 608
rect 1958 542 1961 578
rect 1962 538 1966 541
rect 1982 512 1985 758
rect 1998 752 2001 958
rect 2006 742 2009 1068
rect 2014 962 2017 1208
rect 2022 1152 2025 1268
rect 2030 1192 2033 1268
rect 2054 1222 2057 1258
rect 2062 1242 2065 1408
rect 2042 1218 2046 1221
rect 2070 1202 2073 1458
rect 2078 1422 2081 1428
rect 2086 1402 2089 1508
rect 2098 1498 2102 1501
rect 2078 1352 2081 1388
rect 2086 1372 2089 1378
rect 2094 1352 2097 1428
rect 2110 1422 2113 1528
rect 2102 1372 2105 1408
rect 2078 1242 2081 1318
rect 2062 1152 2065 1158
rect 2070 1152 2073 1198
rect 2086 1182 2089 1348
rect 2098 1328 2102 1331
rect 2094 1312 2097 1318
rect 2094 1262 2097 1268
rect 2024 1103 2026 1107
rect 2030 1103 2033 1107
rect 2038 1103 2040 1107
rect 2046 1082 2049 1098
rect 2022 1022 2025 1028
rect 2022 951 2025 958
rect 2022 948 2030 951
rect 2046 932 2049 998
rect 2014 892 2017 918
rect 2024 903 2026 907
rect 2030 903 2033 907
rect 2038 903 2040 907
rect 2022 822 2025 888
rect 2038 852 2041 868
rect 2046 852 2049 888
rect 2054 872 2057 1148
rect 2070 1122 2073 1138
rect 2078 1132 2081 1138
rect 2062 1092 2065 1108
rect 2070 1052 2073 1078
rect 2062 1032 2065 1048
rect 2066 998 2073 1001
rect 2062 942 2065 948
rect 2034 818 2038 821
rect 2046 772 2049 818
rect 2062 792 2065 918
rect 2070 912 2073 998
rect 2070 842 2073 868
rect 2058 768 2062 771
rect 2018 738 2022 741
rect 2054 732 2057 738
rect 2014 712 2017 728
rect 2024 703 2026 707
rect 2030 703 2033 707
rect 2038 703 2040 707
rect 2014 682 2017 698
rect 2070 682 2073 708
rect 2066 658 2070 661
rect 2078 652 2081 1128
rect 2086 1072 2089 1108
rect 2094 1062 2097 1238
rect 2090 1048 2094 1051
rect 2086 902 2089 928
rect 2086 852 2089 858
rect 2094 772 2097 1048
rect 2102 922 2105 1298
rect 2110 1292 2113 1328
rect 2118 1322 2121 1468
rect 2126 1452 2129 1648
rect 2142 1642 2145 1818
rect 2150 1582 2153 1748
rect 2158 1702 2161 1858
rect 2190 1791 2193 1838
rect 2190 1788 2198 1791
rect 2166 1661 2169 1758
rect 2166 1658 2174 1661
rect 2182 1602 2185 1658
rect 2190 1652 2193 1658
rect 2134 1552 2137 1558
rect 2134 1431 2137 1478
rect 2142 1462 2145 1568
rect 2150 1542 2153 1568
rect 2158 1522 2161 1548
rect 2158 1512 2161 1518
rect 2134 1428 2145 1431
rect 2110 1112 2113 1288
rect 2118 1282 2121 1308
rect 2118 1252 2121 1268
rect 2110 972 2113 1068
rect 2118 1012 2121 1208
rect 2126 1082 2129 1318
rect 2134 1312 2137 1418
rect 2142 1372 2145 1428
rect 2150 1391 2153 1508
rect 2166 1402 2169 1558
rect 2174 1392 2177 1508
rect 2198 1492 2201 1778
rect 2206 1691 2209 1968
rect 2238 1911 2241 1918
rect 2234 1908 2241 1911
rect 2214 1892 2217 1898
rect 2222 1892 2225 1898
rect 2254 1892 2257 2048
rect 2270 1962 2273 2288
rect 2278 1972 2281 2498
rect 2290 2458 2294 2461
rect 2286 2112 2289 2448
rect 2310 2251 2313 2388
rect 2306 2248 2313 2251
rect 2290 2068 2294 2071
rect 2234 1888 2238 1891
rect 2278 1861 2281 1868
rect 2278 1858 2286 1861
rect 2270 1832 2273 1858
rect 2282 1848 2286 1851
rect 2214 1751 2217 1778
rect 2214 1748 2222 1751
rect 2206 1688 2214 1691
rect 2206 1582 2209 1648
rect 2214 1622 2217 1668
rect 2222 1582 2225 1728
rect 2206 1502 2209 1558
rect 2222 1542 2225 1568
rect 2214 1528 2222 1531
rect 2150 1388 2158 1391
rect 2166 1371 2169 1388
rect 2158 1368 2169 1371
rect 2158 1292 2161 1368
rect 2182 1361 2185 1468
rect 2190 1392 2193 1458
rect 2198 1452 2201 1458
rect 2206 1382 2209 1448
rect 2214 1442 2217 1528
rect 2230 1512 2233 1798
rect 2270 1788 2278 1791
rect 2262 1772 2265 1788
rect 2238 1692 2241 1728
rect 2238 1572 2241 1638
rect 2230 1402 2233 1478
rect 2238 1432 2241 1568
rect 2246 1542 2249 1598
rect 2246 1532 2249 1538
rect 2246 1412 2249 1498
rect 2254 1472 2257 1748
rect 2270 1672 2273 1788
rect 2286 1732 2289 1758
rect 2278 1691 2281 1718
rect 2278 1688 2289 1691
rect 2270 1632 2273 1648
rect 2278 1592 2281 1678
rect 2262 1552 2265 1578
rect 2286 1552 2289 1688
rect 2294 1562 2297 2038
rect 2302 1952 2305 2058
rect 2310 2042 2313 2248
rect 2318 2062 2321 2548
rect 2350 2502 2353 2528
rect 2326 2292 2329 2488
rect 2350 2452 2353 2498
rect 2334 2352 2337 2358
rect 2342 2082 2345 2098
rect 2342 2052 2345 2058
rect 2302 1862 2305 1888
rect 2302 1652 2305 1858
rect 2310 1732 2313 1938
rect 2318 1682 2321 1888
rect 2326 1851 2329 1908
rect 2326 1848 2334 1851
rect 2334 1832 2337 1838
rect 2330 1708 2334 1711
rect 2302 1562 2305 1648
rect 2310 1628 2318 1631
rect 2262 1472 2265 1528
rect 2270 1482 2273 1518
rect 2278 1462 2281 1548
rect 2286 1528 2294 1531
rect 2286 1522 2289 1528
rect 2286 1492 2289 1518
rect 2302 1482 2305 1538
rect 2310 1502 2313 1628
rect 2318 1602 2321 1618
rect 2326 1582 2329 1638
rect 2334 1632 2337 1678
rect 2334 1582 2337 1608
rect 2342 1532 2345 1868
rect 2350 1712 2353 2398
rect 2358 2112 2361 2878
rect 2366 2662 2369 2678
rect 2366 2472 2369 2648
rect 2366 2162 2369 2368
rect 2374 1932 2377 2768
rect 2382 2522 2385 3058
rect 2382 2172 2385 2268
rect 2382 2072 2385 2078
rect 2390 2062 2393 2888
rect 2402 2668 2406 2671
rect 2414 2661 2417 2668
rect 2406 2658 2417 2661
rect 2406 2632 2409 2658
rect 2406 2542 2409 2588
rect 2398 2392 2401 2518
rect 2414 2512 2417 2648
rect 2422 2352 2425 2738
rect 2430 2572 2433 2578
rect 2430 2282 2433 2518
rect 2438 2512 2441 2728
rect 2438 2292 2441 2408
rect 2446 2332 2449 3028
rect 2454 2882 2457 3208
rect 2462 2562 2465 3298
rect 2470 3132 2473 3258
rect 2506 3248 2510 3251
rect 2490 3158 2494 3161
rect 2470 3002 2473 3128
rect 2506 3068 2510 3071
rect 2506 3058 2510 3061
rect 2506 2938 2513 2941
rect 2470 2532 2473 2898
rect 2478 2862 2481 2868
rect 2494 2842 2497 2868
rect 2478 2752 2481 2818
rect 2486 2742 2489 2818
rect 2494 2792 2497 2838
rect 2494 2622 2497 2668
rect 2502 2652 2505 2928
rect 2510 2612 2513 2938
rect 2486 2522 2489 2538
rect 2454 2281 2457 2518
rect 2470 2452 2473 2458
rect 2478 2452 2481 2468
rect 2510 2462 2513 2588
rect 2518 2532 2521 3298
rect 2536 3203 2538 3207
rect 2542 3203 2545 3207
rect 2550 3203 2552 3207
rect 2526 2952 2529 3118
rect 2558 3012 2561 3018
rect 2536 3003 2538 3007
rect 2542 3003 2545 3007
rect 2550 3003 2552 3007
rect 2562 2858 2566 2861
rect 2574 2852 2577 3268
rect 2578 2848 2585 2851
rect 2582 2822 2585 2848
rect 2590 2811 2593 3048
rect 2582 2808 2593 2811
rect 2536 2803 2538 2807
rect 2542 2803 2545 2807
rect 2550 2803 2552 2807
rect 2554 2758 2558 2761
rect 2526 2562 2529 2718
rect 2536 2603 2538 2607
rect 2542 2603 2545 2607
rect 2550 2603 2552 2607
rect 2558 2582 2561 2598
rect 2530 2528 2534 2531
rect 2546 2458 2550 2461
rect 2454 2278 2462 2281
rect 2398 2052 2401 2078
rect 2382 1922 2385 1948
rect 2358 1702 2361 1728
rect 2350 1692 2353 1698
rect 2374 1691 2377 1728
rect 2358 1688 2377 1691
rect 2270 1452 2273 1458
rect 2302 1442 2305 1458
rect 2182 1358 2190 1361
rect 2182 1332 2185 1348
rect 2166 1302 2169 1318
rect 2134 1268 2142 1271
rect 2134 1202 2137 1268
rect 2142 1232 2145 1248
rect 2142 1152 2145 1158
rect 2134 1062 2137 1108
rect 2150 1092 2153 1268
rect 2158 1081 2161 1258
rect 2166 1092 2169 1268
rect 2174 1182 2177 1288
rect 2182 1282 2185 1298
rect 2182 1172 2185 1248
rect 2198 1242 2201 1358
rect 2206 1292 2209 1378
rect 2222 1362 2225 1378
rect 2230 1372 2233 1388
rect 2238 1372 2241 1398
rect 2214 1332 2217 1348
rect 2206 1232 2209 1238
rect 2190 1228 2198 1231
rect 2190 1212 2193 1228
rect 2174 1142 2177 1148
rect 2150 1078 2161 1081
rect 2150 1032 2153 1078
rect 2162 1058 2166 1061
rect 2174 1042 2177 1088
rect 2190 1042 2193 1068
rect 2178 958 2182 961
rect 2102 892 2105 898
rect 2118 872 2121 958
rect 2158 902 2161 948
rect 2086 662 2089 678
rect 2110 672 2113 768
rect 2118 732 2121 768
rect 2134 752 2137 898
rect 2150 812 2153 868
rect 2142 762 2145 798
rect 2158 762 2161 838
rect 2158 722 2161 738
rect 1990 552 1993 578
rect 1934 412 1937 508
rect 1942 401 1945 408
rect 1934 398 1945 401
rect 1934 212 1937 398
rect 1962 368 1966 371
rect 1942 312 1945 358
rect 1990 272 1993 548
rect 1998 342 2001 648
rect 2082 638 2089 641
rect 2086 602 2089 638
rect 2024 503 2026 507
rect 2030 503 2033 507
rect 2038 503 2040 507
rect 2110 472 2113 668
rect 2126 642 2129 678
rect 2150 662 2153 668
rect 2134 542 2137 658
rect 2166 612 2169 938
rect 2174 752 2177 888
rect 2182 812 2185 948
rect 2174 482 2177 698
rect 2182 482 2185 788
rect 2170 478 2174 481
rect 2006 468 2014 471
rect 2006 442 2009 468
rect 2174 452 2177 468
rect 2102 352 2105 398
rect 2114 328 2118 331
rect 2006 312 2009 328
rect 2014 302 2017 318
rect 2024 303 2026 307
rect 2030 303 2033 307
rect 2038 303 2040 307
rect 1974 242 1977 268
rect 1990 242 1993 268
rect 1982 232 1985 238
rect 1798 142 1801 148
rect 1806 142 1809 148
rect 1966 142 1969 228
rect 1710 112 1713 128
rect 1798 122 1801 128
rect 1798 82 1801 98
rect 1618 58 1622 61
rect 1630 52 1633 58
rect 1806 52 1809 118
rect 1886 81 1889 98
rect 1882 78 1889 81
rect 1922 78 1926 81
rect 1970 78 1974 81
rect 1982 81 1985 178
rect 2046 162 2049 328
rect 2066 268 2070 271
rect 2086 252 2089 258
rect 2098 158 2102 161
rect 2062 132 2065 158
rect 2024 103 2026 107
rect 2030 103 2033 107
rect 2038 103 2040 107
rect 2118 102 2121 158
rect 2126 132 2129 338
rect 2158 282 2161 308
rect 2190 272 2193 968
rect 2198 942 2201 1168
rect 2222 1102 2225 1328
rect 2230 1242 2233 1318
rect 2246 1312 2249 1318
rect 2246 1272 2249 1288
rect 2206 1072 2209 1078
rect 2206 962 2209 998
rect 2214 932 2217 1078
rect 2230 1072 2233 1128
rect 2222 1032 2225 1038
rect 2238 992 2241 1158
rect 2254 1152 2257 1368
rect 2270 1352 2273 1358
rect 2262 1262 2265 1348
rect 2262 1102 2265 1258
rect 2270 1242 2273 1338
rect 2258 1088 2262 1091
rect 2246 1082 2249 1088
rect 2230 968 2238 971
rect 2230 962 2233 968
rect 2206 871 2209 878
rect 2202 868 2209 871
rect 2230 851 2233 908
rect 2242 868 2246 871
rect 2230 848 2238 851
rect 2198 732 2201 748
rect 2206 672 2209 808
rect 2230 742 2233 768
rect 2254 632 2257 1048
rect 2262 1002 2265 1068
rect 2270 1012 2273 1168
rect 2278 1011 2281 1358
rect 2286 1282 2289 1288
rect 2286 1232 2289 1258
rect 2294 1142 2297 1388
rect 2302 1302 2305 1328
rect 2302 1232 2305 1238
rect 2310 1162 2313 1338
rect 2310 1122 2313 1128
rect 2294 1052 2297 1088
rect 2294 1012 2297 1048
rect 2278 1008 2286 1011
rect 2270 991 2273 998
rect 2262 988 2273 991
rect 2262 972 2265 988
rect 2278 892 2281 978
rect 2262 872 2265 888
rect 2286 822 2289 978
rect 2302 942 2305 1048
rect 2310 922 2313 1078
rect 2310 872 2313 878
rect 2282 748 2286 751
rect 2274 738 2278 741
rect 2294 722 2297 838
rect 2278 718 2286 721
rect 2138 268 2142 271
rect 2142 152 2145 158
rect 2142 112 2145 128
rect 2166 112 2169 238
rect 2174 122 2177 178
rect 2182 152 2185 158
rect 1982 78 1990 81
rect 2014 81 2017 98
rect 2010 78 2017 81
rect 2058 78 2062 81
rect 1902 52 1905 78
rect 2006 62 2009 68
rect 2198 62 2201 508
rect 2214 322 2217 358
rect 2238 251 2241 258
rect 2234 248 2241 251
rect 2222 62 2225 68
rect 2238 62 2241 118
rect 2246 112 2249 418
rect 2278 402 2281 718
rect 2302 622 2305 868
rect 2318 732 2321 1528
rect 2334 1492 2337 1498
rect 2334 1462 2337 1478
rect 2342 1252 2345 1488
rect 2350 1382 2353 1678
rect 2358 1622 2361 1688
rect 2366 1622 2369 1628
rect 2358 1592 2361 1598
rect 2358 1562 2361 1568
rect 2366 1552 2369 1588
rect 2358 1492 2361 1498
rect 2358 1432 2361 1468
rect 2366 1442 2369 1478
rect 2350 1362 2353 1378
rect 2358 1332 2361 1398
rect 2366 1362 2369 1368
rect 2350 1282 2353 1308
rect 2358 1271 2361 1278
rect 2350 1268 2361 1271
rect 2334 1212 2337 1228
rect 2350 1222 2353 1268
rect 2326 1032 2329 1058
rect 2334 941 2337 1208
rect 2350 1132 2353 1208
rect 2350 1082 2353 1118
rect 2330 938 2337 941
rect 2342 901 2345 1008
rect 2350 952 2353 968
rect 2342 898 2350 901
rect 2334 762 2337 768
rect 2302 452 2305 468
rect 2310 452 2313 678
rect 2270 202 2273 328
rect 2318 292 2321 688
rect 2342 662 2345 708
rect 2358 582 2361 1218
rect 2366 1092 2369 1328
rect 2374 1302 2377 1678
rect 2382 1572 2385 1868
rect 2406 1862 2409 2248
rect 2470 2162 2473 2358
rect 2478 2272 2481 2448
rect 2486 2272 2489 2348
rect 2506 2328 2510 2331
rect 2418 2078 2422 2081
rect 2418 2048 2422 2051
rect 2430 1882 2433 1998
rect 2438 1932 2441 2008
rect 2446 2002 2449 2078
rect 2422 1762 2425 1808
rect 2406 1732 2409 1748
rect 2398 1681 2401 1718
rect 2394 1678 2401 1681
rect 2406 1622 2409 1678
rect 2422 1652 2425 1728
rect 2430 1722 2433 1758
rect 2438 1632 2441 1818
rect 2422 1582 2425 1628
rect 2446 1561 2449 1998
rect 2478 1952 2481 2098
rect 2486 2062 2489 2268
rect 2518 2252 2521 2438
rect 2526 2422 2529 2428
rect 2536 2403 2538 2407
rect 2542 2403 2545 2407
rect 2550 2403 2552 2407
rect 2558 2332 2561 2578
rect 2574 2282 2577 2798
rect 2582 2492 2585 2808
rect 2590 2712 2593 2798
rect 2590 2662 2593 2668
rect 2590 2562 2593 2608
rect 2590 2462 2593 2538
rect 2598 2492 2601 2868
rect 2606 2582 2609 2878
rect 2630 2672 2633 3298
rect 2638 2652 2641 2748
rect 2646 2642 2649 3298
rect 2762 3258 2766 3261
rect 2678 3142 2681 3258
rect 2706 3158 2710 3161
rect 2770 3138 2774 3141
rect 2654 2622 2657 2698
rect 2618 2578 2622 2581
rect 2594 2358 2601 2361
rect 2582 2332 2585 2358
rect 2598 2342 2601 2358
rect 2598 2322 2601 2338
rect 2494 2238 2502 2241
rect 2494 2142 2497 2238
rect 2566 2232 2569 2238
rect 2514 2208 2518 2211
rect 2536 2203 2538 2207
rect 2542 2203 2545 2207
rect 2550 2203 2552 2207
rect 2530 2138 2534 2141
rect 2526 2122 2529 2138
rect 2574 2132 2577 2278
rect 2582 2112 2585 2278
rect 2598 2272 2601 2278
rect 2486 2042 2489 2048
rect 2478 1902 2481 1928
rect 2486 1902 2489 1908
rect 2486 1842 2489 1888
rect 2454 1751 2457 1768
rect 2454 1748 2462 1751
rect 2454 1682 2457 1738
rect 2438 1558 2449 1561
rect 2454 1562 2457 1648
rect 2462 1592 2465 1708
rect 2470 1662 2473 1788
rect 2486 1732 2489 1808
rect 2382 1452 2385 1538
rect 2390 1512 2393 1548
rect 2398 1522 2401 1538
rect 2422 1512 2425 1558
rect 2390 1432 2393 1508
rect 2418 1448 2422 1451
rect 2382 1342 2385 1418
rect 2390 1372 2393 1428
rect 2406 1392 2409 1408
rect 2406 1351 2409 1378
rect 2402 1348 2409 1351
rect 2374 1272 2377 1288
rect 2382 1281 2385 1338
rect 2382 1278 2390 1281
rect 2386 1268 2390 1271
rect 2366 952 2369 1078
rect 2374 942 2377 1268
rect 2398 1242 2401 1308
rect 2406 1282 2409 1298
rect 2414 1242 2417 1278
rect 2422 1222 2425 1428
rect 2430 1272 2433 1348
rect 2438 1272 2441 1558
rect 2450 1548 2457 1551
rect 2454 1542 2457 1548
rect 2478 1502 2481 1618
rect 2478 1472 2481 1498
rect 2446 1402 2449 1448
rect 2454 1312 2457 1448
rect 2470 1392 2473 1408
rect 2478 1382 2481 1438
rect 2462 1291 2465 1368
rect 2470 1322 2473 1328
rect 2474 1308 2481 1311
rect 2458 1288 2465 1291
rect 2442 1258 2446 1261
rect 2430 1202 2433 1238
rect 2382 1152 2385 1178
rect 2478 1162 2481 1308
rect 2486 1222 2489 1598
rect 2494 1482 2497 1798
rect 2502 1761 2505 1938
rect 2510 1802 2513 2008
rect 2526 1942 2529 2008
rect 2536 2003 2538 2007
rect 2542 2003 2545 2007
rect 2550 2003 2552 2007
rect 2536 1803 2538 1807
rect 2542 1803 2545 1807
rect 2550 1803 2552 1807
rect 2558 1802 2561 1818
rect 2502 1758 2513 1761
rect 2510 1702 2513 1758
rect 2522 1748 2526 1751
rect 2550 1702 2553 1778
rect 2546 1688 2550 1691
rect 2510 1582 2513 1688
rect 2558 1682 2561 1688
rect 2522 1658 2526 1661
rect 2526 1632 2529 1658
rect 2534 1622 2537 1658
rect 2566 1632 2569 1978
rect 2574 1752 2577 1818
rect 2582 1811 2585 1848
rect 2590 1822 2593 2038
rect 2606 1952 2609 2538
rect 2622 2442 2625 2488
rect 2638 2302 2641 2408
rect 2646 2302 2649 2398
rect 2670 2302 2673 2328
rect 2678 2322 2681 3138
rect 2782 3062 2785 3148
rect 2638 2022 2641 2248
rect 2646 2142 2649 2298
rect 2582 1808 2593 1811
rect 2574 1662 2577 1718
rect 2536 1603 2538 1607
rect 2542 1603 2545 1607
rect 2550 1603 2552 1607
rect 2582 1602 2585 1798
rect 2590 1752 2593 1808
rect 2606 1752 2609 1788
rect 2590 1692 2593 1748
rect 2614 1722 2617 1828
rect 2614 1682 2617 1698
rect 2526 1592 2529 1598
rect 2590 1572 2593 1648
rect 2602 1638 2609 1641
rect 2502 1562 2505 1568
rect 2598 1562 2601 1628
rect 2554 1548 2561 1551
rect 2558 1542 2561 1548
rect 2538 1528 2542 1531
rect 2502 1362 2505 1398
rect 2382 1071 2385 1148
rect 2478 1142 2481 1148
rect 2406 1122 2409 1138
rect 2382 1068 2393 1071
rect 2390 952 2393 1068
rect 2390 932 2393 948
rect 2366 652 2369 718
rect 2390 702 2393 798
rect 2398 692 2401 1088
rect 2414 1072 2417 1078
rect 2430 1002 2433 1078
rect 2438 1072 2441 1088
rect 2430 991 2433 998
rect 2426 988 2433 991
rect 2446 872 2449 988
rect 2478 892 2481 1128
rect 2486 1002 2489 1168
rect 2494 1042 2497 1318
rect 2466 878 2470 881
rect 2410 858 2417 861
rect 2414 852 2417 858
rect 2414 761 2417 778
rect 2410 758 2417 761
rect 2418 728 2425 731
rect 2414 681 2417 688
rect 2410 678 2417 681
rect 2374 662 2377 668
rect 2422 582 2425 728
rect 2430 672 2433 858
rect 2438 672 2441 788
rect 2330 478 2334 481
rect 2314 268 2318 271
rect 2326 268 2334 271
rect 2262 62 2265 118
rect 2282 98 2289 101
rect 2286 92 2289 98
rect 2234 58 2238 61
rect 1802 48 1806 51
rect 2294 42 2297 258
rect 2302 182 2305 248
rect 2326 222 2329 268
rect 2326 132 2329 218
rect 2330 108 2334 111
rect 2318 102 2321 108
rect 2326 92 2329 98
rect 2334 62 2337 78
rect 2342 12 2345 478
rect 2370 438 2377 441
rect 2358 332 2361 348
rect 2374 242 2377 438
rect 2382 272 2385 498
rect 2446 482 2449 818
rect 2502 802 2505 1348
rect 2510 1342 2513 1518
rect 2558 1472 2561 1528
rect 2566 1522 2569 1548
rect 2574 1522 2577 1538
rect 2566 1482 2569 1518
rect 2582 1472 2585 1558
rect 2550 1462 2553 1468
rect 2546 1448 2550 1451
rect 2510 1292 2513 1318
rect 2518 1292 2521 1368
rect 2526 1362 2529 1438
rect 2536 1403 2538 1407
rect 2542 1403 2545 1407
rect 2550 1403 2552 1407
rect 2526 1332 2529 1338
rect 2526 1312 2529 1328
rect 2510 1092 2513 1258
rect 2536 1203 2538 1207
rect 2542 1203 2545 1207
rect 2550 1203 2552 1207
rect 2518 1141 2521 1148
rect 2518 1138 2526 1141
rect 2522 1128 2529 1131
rect 2546 1128 2550 1131
rect 2518 1012 2521 1028
rect 2526 1022 2529 1128
rect 2558 1082 2561 1458
rect 2550 1042 2553 1068
rect 2536 1003 2538 1007
rect 2542 1003 2545 1007
rect 2550 1003 2552 1007
rect 2466 738 2470 741
rect 2482 728 2486 731
rect 2498 638 2502 641
rect 2390 262 2393 458
rect 2422 322 2425 468
rect 2470 401 2473 418
rect 2470 398 2478 401
rect 2470 382 2473 398
rect 2438 312 2441 348
rect 2462 312 2465 338
rect 2398 272 2401 278
rect 2382 211 2385 258
rect 2378 208 2385 211
rect 2462 192 2465 308
rect 2510 292 2513 868
rect 2518 522 2521 868
rect 2536 803 2538 807
rect 2542 803 2545 807
rect 2550 803 2552 807
rect 2526 742 2529 798
rect 2526 612 2529 678
rect 2536 603 2538 607
rect 2542 603 2545 607
rect 2550 603 2552 607
rect 2536 403 2538 407
rect 2542 403 2545 407
rect 2550 403 2552 407
rect 2558 302 2561 1048
rect 2566 912 2569 1448
rect 2590 1412 2593 1548
rect 2598 1462 2601 1548
rect 2574 1052 2577 1388
rect 2582 1352 2585 1388
rect 2598 1361 2601 1378
rect 2594 1358 2601 1361
rect 2582 982 2585 1338
rect 2590 1292 2593 1328
rect 2598 1302 2601 1328
rect 2598 982 2601 1218
rect 2606 1192 2609 1638
rect 2614 1352 2617 1668
rect 2614 1152 2617 1288
rect 2622 1172 2625 1898
rect 2630 1722 2633 1868
rect 2630 1492 2633 1658
rect 2638 1622 2641 2018
rect 2646 1832 2649 2138
rect 2654 2032 2657 2048
rect 2654 1792 2657 2018
rect 2662 1881 2665 2238
rect 2678 2002 2681 2188
rect 2686 2172 2689 2368
rect 2702 2352 2705 2748
rect 2694 1982 2697 2318
rect 2678 1958 2686 1961
rect 2678 1952 2681 1958
rect 2702 1942 2705 2348
rect 2718 2061 2721 2718
rect 2734 2672 2737 2758
rect 2742 2642 2745 2838
rect 2766 2692 2769 3038
rect 2762 2668 2766 2671
rect 2774 2662 2777 2898
rect 2710 2058 2721 2061
rect 2710 1912 2713 2058
rect 2662 1878 2678 1881
rect 2658 1788 2662 1791
rect 2646 1602 2649 1788
rect 2654 1662 2657 1768
rect 2670 1742 2673 1878
rect 2686 1872 2689 1878
rect 2702 1868 2710 1871
rect 2678 1792 2681 1808
rect 2678 1692 2681 1708
rect 2686 1692 2689 1698
rect 2654 1632 2657 1658
rect 2662 1652 2665 1658
rect 2630 1272 2633 1408
rect 2638 1352 2641 1548
rect 2646 1532 2649 1568
rect 2658 1558 2662 1561
rect 2662 1492 2665 1508
rect 2654 1342 2657 1348
rect 2642 1268 2646 1271
rect 2630 1252 2633 1258
rect 2638 1202 2641 1268
rect 2654 1242 2657 1318
rect 2670 1312 2673 1488
rect 2678 1472 2681 1478
rect 2678 1372 2681 1468
rect 2686 1462 2689 1608
rect 2694 1402 2697 1758
rect 2702 1752 2705 1868
rect 2718 1822 2721 2048
rect 2726 1912 2729 2488
rect 2742 2112 2745 2418
rect 2766 2372 2769 2638
rect 2774 2442 2777 2548
rect 2782 2462 2785 3058
rect 2790 2872 2793 3288
rect 2790 2742 2793 2868
rect 2806 2852 2809 3298
rect 2854 3082 2857 3268
rect 2878 2942 2881 2958
rect 2790 2632 2793 2738
rect 2798 2562 2801 2728
rect 2806 2681 2809 2828
rect 2814 2692 2817 2758
rect 2806 2678 2817 2681
rect 2746 2068 2750 2071
rect 2734 1992 2737 2028
rect 2750 1972 2753 1988
rect 2742 1921 2745 1968
rect 2738 1918 2745 1921
rect 2758 1912 2761 2308
rect 2766 1992 2769 2208
rect 2774 2072 2777 2338
rect 2782 2062 2785 2458
rect 2798 2202 2801 2528
rect 2806 2222 2809 2338
rect 2686 1332 2689 1358
rect 2702 1342 2705 1718
rect 2718 1681 2721 1738
rect 2714 1678 2721 1681
rect 2710 1382 2713 1598
rect 2694 1332 2697 1338
rect 2614 1082 2617 1148
rect 2606 972 2609 978
rect 2566 782 2569 798
rect 2566 442 2569 708
rect 2574 532 2577 928
rect 2638 912 2641 1188
rect 2598 692 2601 788
rect 2614 582 2617 888
rect 2634 778 2638 781
rect 2626 728 2630 731
rect 2646 662 2649 1178
rect 2654 952 2657 1068
rect 2662 942 2665 1118
rect 2670 902 2673 1308
rect 2686 862 2689 1258
rect 2702 1252 2705 1318
rect 2710 1252 2713 1378
rect 2718 1262 2721 1618
rect 2726 1612 2729 1858
rect 2758 1791 2761 1848
rect 2766 1802 2769 1948
rect 2758 1788 2769 1791
rect 2734 1651 2737 1708
rect 2734 1648 2742 1651
rect 2758 1612 2761 1678
rect 2742 1572 2745 1578
rect 2754 1558 2758 1561
rect 2754 1528 2758 1531
rect 2734 1522 2737 1528
rect 2726 1512 2729 1518
rect 2726 1242 2729 1388
rect 2734 1302 2737 1498
rect 2758 1472 2761 1478
rect 2742 1452 2745 1468
rect 2742 1362 2745 1368
rect 2742 1332 2745 1338
rect 2742 1242 2745 1258
rect 2750 1172 2753 1418
rect 2758 1362 2761 1468
rect 2766 1452 2769 1788
rect 2774 1572 2777 1658
rect 2758 1312 2761 1338
rect 2766 1332 2769 1448
rect 2774 1321 2777 1568
rect 2766 1318 2777 1321
rect 2710 1141 2713 1148
rect 2706 1138 2713 1141
rect 2738 1138 2745 1141
rect 2718 1102 2721 1128
rect 2742 1122 2745 1138
rect 2758 1112 2761 1168
rect 2766 1082 2769 1318
rect 2774 1242 2777 1248
rect 2774 1112 2777 1238
rect 2782 1162 2785 2058
rect 2794 2038 2798 2041
rect 2814 1982 2817 2678
rect 2822 2582 2825 2668
rect 2838 2661 2841 2738
rect 2834 2658 2841 2661
rect 2858 2658 2865 2661
rect 2838 2482 2841 2638
rect 2850 2538 2854 2541
rect 2790 1502 2793 1778
rect 2798 1662 2801 1758
rect 2806 1702 2809 1738
rect 2814 1642 2817 1748
rect 2822 1602 2825 2278
rect 2830 2122 2833 2468
rect 2854 2382 2857 2398
rect 2854 2252 2857 2378
rect 2862 2342 2865 2658
rect 2870 2552 2873 2578
rect 2878 2421 2881 2938
rect 2886 2732 2889 2738
rect 2910 2702 2913 3058
rect 2918 2682 2921 3258
rect 2926 2772 2929 3288
rect 3002 3138 3009 3141
rect 2934 2932 2937 2938
rect 2934 2722 2937 2928
rect 2950 2718 2958 2721
rect 2918 2502 2921 2678
rect 2938 2608 2945 2611
rect 2942 2592 2945 2608
rect 2950 2562 2953 2718
rect 2990 2682 2993 2998
rect 3006 2992 3009 3138
rect 3040 3103 3042 3107
rect 3046 3103 3049 3107
rect 3054 3103 3056 3107
rect 3086 3052 3089 3298
rect 3506 3278 3510 3281
rect 3298 3268 3302 3271
rect 3514 3268 3518 3271
rect 3122 3258 3126 3261
rect 3094 3252 3097 3258
rect 3102 3162 3105 3178
rect 3174 3112 3177 3258
rect 3122 2918 3129 2921
rect 3040 2903 3042 2907
rect 3046 2903 3049 2907
rect 3054 2903 3056 2907
rect 3126 2892 3129 2918
rect 2998 2862 3001 2868
rect 2878 2418 2886 2421
rect 2866 2248 2870 2251
rect 2874 2028 2878 2031
rect 2886 2012 2889 2418
rect 2894 2002 2897 2318
rect 2902 2101 2905 2308
rect 2918 2302 2921 2418
rect 2950 2362 2953 2488
rect 2958 2462 2961 2478
rect 2910 2112 2913 2158
rect 2902 2098 2913 2101
rect 2902 2052 2905 2058
rect 2866 1988 2870 1991
rect 2842 1878 2846 1881
rect 2842 1858 2846 1861
rect 2830 1722 2833 1768
rect 2854 1572 2857 1898
rect 2842 1548 2846 1551
rect 2802 1528 2806 1531
rect 2818 1528 2825 1531
rect 2710 922 2713 1058
rect 2718 912 2721 1068
rect 2658 728 2665 731
rect 2662 712 2665 728
rect 2502 272 2505 278
rect 2490 268 2494 271
rect 2478 242 2481 258
rect 2558 252 2561 278
rect 2566 252 2569 438
rect 2574 352 2577 528
rect 2638 492 2641 568
rect 2670 542 2673 838
rect 2678 822 2681 858
rect 2706 838 2710 841
rect 2706 818 2710 821
rect 2678 542 2681 818
rect 2726 742 2729 1078
rect 2742 771 2745 828
rect 2738 768 2745 771
rect 2750 742 2753 748
rect 2686 648 2694 651
rect 2662 522 2665 538
rect 2686 522 2689 648
rect 2674 518 2681 521
rect 2638 482 2641 488
rect 2602 468 2606 471
rect 2586 348 2590 351
rect 2486 212 2489 248
rect 2350 152 2353 158
rect 2366 142 2369 148
rect 2362 108 2366 111
rect 2362 58 2366 61
rect 2374 12 2377 178
rect 2398 132 2401 138
rect 2406 132 2409 138
rect 2406 102 2409 118
rect 2390 61 2393 68
rect 2386 58 2393 61
rect 2414 11 2417 148
rect 2478 102 2481 128
rect 2486 122 2489 168
rect 2502 92 2505 128
rect 2526 112 2529 218
rect 2536 203 2538 207
rect 2542 203 2545 207
rect 2550 203 2552 207
rect 2462 52 2465 58
rect 2574 32 2577 308
rect 2582 292 2585 338
rect 2678 322 2681 518
rect 2690 448 2694 451
rect 2694 372 2697 448
rect 2702 362 2705 508
rect 2710 312 2713 618
rect 2734 482 2737 488
rect 2742 452 2745 658
rect 2614 272 2617 298
rect 2690 258 2694 261
rect 2710 232 2713 298
rect 2718 232 2721 238
rect 2666 158 2670 161
rect 2582 82 2585 88
rect 2590 42 2593 128
rect 2678 21 2681 158
rect 2750 142 2753 148
rect 2710 92 2713 108
rect 2686 42 2689 78
rect 2750 62 2753 78
rect 2678 18 2686 21
rect 2758 12 2761 748
rect 2766 742 2769 958
rect 2774 512 2777 1098
rect 2766 321 2769 498
rect 2766 318 2774 321
rect 2766 308 2774 311
rect 2766 222 2769 308
rect 2770 138 2774 141
rect 2782 62 2785 1158
rect 2790 662 2793 1438
rect 2798 1332 2801 1438
rect 2822 1422 2825 1528
rect 2854 1512 2857 1548
rect 2830 1382 2833 1388
rect 2830 1352 2833 1358
rect 2854 1352 2857 1508
rect 2862 1392 2865 1588
rect 2870 1552 2873 1978
rect 2878 1662 2881 1978
rect 2910 1942 2913 2098
rect 2918 2022 2921 2108
rect 2926 1992 2929 2338
rect 2934 2152 2937 2158
rect 2942 2142 2945 2358
rect 2942 2082 2945 2138
rect 2918 1952 2921 1958
rect 2926 1952 2929 1958
rect 2942 1941 2945 1948
rect 2938 1938 2945 1941
rect 2950 1932 2953 2328
rect 2958 2162 2961 2448
rect 2974 2362 2977 2568
rect 2990 2472 2993 2658
rect 2998 2632 3001 2858
rect 3018 2768 3022 2771
rect 3030 2692 3033 2718
rect 3040 2703 3042 2707
rect 3046 2703 3049 2707
rect 3054 2703 3056 2707
rect 3040 2503 3042 2507
rect 3046 2503 3049 2507
rect 3054 2503 3056 2507
rect 3126 2341 3129 2488
rect 3134 2392 3137 2838
rect 3150 2512 3153 2868
rect 3166 2758 3174 2761
rect 3166 2732 3169 2758
rect 3182 2662 3185 2768
rect 3198 2762 3201 2888
rect 3182 2582 3185 2658
rect 3142 2442 3145 2448
rect 3122 2338 3129 2341
rect 3142 2342 3145 2438
rect 3158 2432 3161 2538
rect 3166 2472 3169 2508
rect 3174 2472 3177 2478
rect 2966 2162 2969 2318
rect 2974 1992 2977 2318
rect 3040 2303 3042 2307
rect 3046 2303 3049 2307
rect 3054 2303 3056 2307
rect 3106 2288 3110 2291
rect 3090 2248 3094 2251
rect 2990 2222 2993 2228
rect 2998 2172 3001 2218
rect 3030 2102 3033 2128
rect 3040 2103 3042 2107
rect 3046 2103 3049 2107
rect 3054 2103 3056 2107
rect 3134 2082 3137 2288
rect 3150 2272 3153 2278
rect 3190 2222 3193 2448
rect 3198 2291 3201 2358
rect 3206 2352 3209 2958
rect 3198 2288 3206 2291
rect 3202 2268 3206 2271
rect 3154 2148 3158 2151
rect 3190 2148 3198 2151
rect 3150 2062 3153 2068
rect 3042 2048 3046 2051
rect 3010 2038 3014 2041
rect 3010 1968 3014 1971
rect 3058 1938 3062 1941
rect 2910 1908 2918 1911
rect 2910 1832 2913 1908
rect 2910 1671 2913 1728
rect 2906 1668 2913 1671
rect 2918 1642 2921 1878
rect 2882 1628 2886 1631
rect 2878 1482 2881 1628
rect 2890 1558 2894 1561
rect 2898 1548 2902 1551
rect 2894 1472 2897 1528
rect 2806 1332 2809 1338
rect 2814 1262 2817 1328
rect 2854 1322 2857 1348
rect 2834 1298 2838 1301
rect 2846 1292 2849 1318
rect 2854 1292 2857 1298
rect 2838 1252 2841 1278
rect 2862 1272 2865 1388
rect 2874 1298 2878 1301
rect 2830 1238 2838 1241
rect 2798 542 2801 548
rect 2794 478 2798 481
rect 2790 442 2793 468
rect 2790 152 2793 438
rect 2798 272 2801 448
rect 2806 282 2809 1228
rect 2814 1082 2817 1098
rect 2814 472 2817 528
rect 2814 442 2817 468
rect 2830 432 2833 1238
rect 2878 1142 2881 1268
rect 2886 1172 2889 1448
rect 2894 1412 2897 1458
rect 2902 1432 2905 1478
rect 2910 1422 2913 1558
rect 2926 1532 2929 1818
rect 2934 1792 2937 1818
rect 2942 1722 2945 1748
rect 2938 1678 2942 1681
rect 2922 1508 2926 1511
rect 2926 1462 2929 1468
rect 2902 1262 2905 1378
rect 2918 1332 2921 1338
rect 2926 1322 2929 1328
rect 2838 692 2841 748
rect 2846 552 2849 1138
rect 2862 1122 2865 1128
rect 2910 1082 2913 1298
rect 2922 1278 2926 1281
rect 2934 1272 2937 1528
rect 2922 1258 2926 1261
rect 2942 1261 2945 1568
rect 2950 1472 2953 1928
rect 2934 1258 2945 1261
rect 2858 1048 2862 1051
rect 2894 932 2897 968
rect 2822 342 2825 368
rect 2798 252 2801 268
rect 2818 258 2822 261
rect 2842 158 2846 161
rect 2826 148 2830 151
rect 2810 128 2814 131
rect 2798 82 2801 88
rect 2854 81 2857 878
rect 2862 581 2865 888
rect 2870 722 2873 858
rect 2894 711 2897 908
rect 2902 852 2905 858
rect 2902 752 2905 778
rect 2890 708 2897 711
rect 2910 702 2913 1078
rect 2918 1052 2921 1058
rect 2918 972 2921 1028
rect 2926 982 2929 1068
rect 2934 922 2937 1258
rect 2950 1182 2953 1348
rect 2958 1172 2961 1938
rect 3040 1903 3042 1907
rect 3046 1903 3049 1907
rect 3054 1903 3056 1907
rect 2966 1452 2969 1868
rect 2974 1692 2977 1898
rect 3002 1868 3006 1871
rect 3002 1858 3006 1861
rect 3002 1758 3006 1761
rect 2982 1752 2985 1758
rect 2982 1681 2985 1688
rect 2978 1678 2985 1681
rect 2966 1202 2969 1448
rect 2974 1402 2977 1588
rect 2974 1322 2977 1328
rect 2982 1302 2985 1468
rect 2990 1312 2993 1418
rect 2998 1351 3001 1498
rect 2998 1348 3006 1351
rect 2978 1278 2982 1281
rect 2978 1268 2982 1271
rect 2962 1138 2966 1141
rect 2890 658 2894 661
rect 2862 578 2870 581
rect 2878 352 2881 368
rect 2902 232 2905 448
rect 2846 78 2857 81
rect 2766 12 2769 18
rect 2846 12 2849 78
rect 2862 72 2865 168
rect 2926 162 2929 838
rect 2942 542 2945 1068
rect 2974 1022 2977 1258
rect 2982 1152 2985 1158
rect 2954 1008 2958 1011
rect 2966 892 2969 978
rect 2982 882 2985 948
rect 2970 738 2974 741
rect 2942 352 2945 398
rect 2938 338 2942 341
rect 2950 162 2953 428
rect 2870 152 2873 158
rect 2874 128 2878 131
rect 2886 122 2889 148
rect 2886 82 2889 108
rect 2894 92 2897 148
rect 2902 122 2905 158
rect 2934 142 2937 158
rect 2942 142 2945 148
rect 2958 102 2961 728
rect 2990 692 2993 1278
rect 2998 1092 3001 1328
rect 2998 742 3001 948
rect 2974 322 2977 338
rect 2978 308 2985 311
rect 2982 202 2985 308
rect 2990 222 2993 448
rect 3006 282 3009 1328
rect 3014 542 3017 1858
rect 3030 1692 3033 1708
rect 3040 1703 3042 1707
rect 3046 1703 3049 1707
rect 3054 1703 3056 1707
rect 3034 1678 3038 1681
rect 3062 1592 3065 1888
rect 3078 1872 3081 1888
rect 3070 1752 3073 1798
rect 3078 1622 3081 1868
rect 3118 1852 3121 2008
rect 3126 1892 3129 2038
rect 3126 1862 3129 1868
rect 3154 1848 3161 1851
rect 3146 1818 3153 1821
rect 3086 1572 3089 1758
rect 3150 1742 3153 1818
rect 3158 1802 3161 1848
rect 3166 1692 3169 1838
rect 3190 1792 3193 2148
rect 3198 2072 3201 2078
rect 3198 1952 3201 1958
rect 3202 1938 3206 1941
rect 3214 1912 3217 3188
rect 3298 3158 3302 3161
rect 3274 2958 3278 2961
rect 3266 2928 3270 2931
rect 3230 2682 3233 2748
rect 3254 2652 3257 2748
rect 3262 2672 3265 2848
rect 3222 2152 3225 2618
rect 3242 2528 3246 2531
rect 3254 2462 3257 2648
rect 3270 2432 3273 2658
rect 3274 2428 3281 2431
rect 3278 2322 3281 2428
rect 3234 2248 3238 2251
rect 3242 2238 3246 2241
rect 3242 2218 3246 2221
rect 3286 2131 3289 2718
rect 3294 2232 3297 2238
rect 3286 2128 3294 2131
rect 3302 2121 3305 3108
rect 3310 3012 3313 3268
rect 3322 3148 3326 3151
rect 3310 2592 3313 3008
rect 3334 2878 3342 2881
rect 3318 2822 3321 2878
rect 3334 2842 3337 2878
rect 3318 2642 3321 2728
rect 3334 2482 3337 2668
rect 3314 2328 3318 2331
rect 3322 2288 3326 2291
rect 3294 2118 3305 2121
rect 3238 2072 3241 2108
rect 3262 1962 3265 2108
rect 3270 1952 3273 1958
rect 3174 1691 3177 1718
rect 3174 1688 3182 1691
rect 3182 1652 3185 1668
rect 3078 1561 3081 1568
rect 3074 1558 3081 1561
rect 3040 1503 3042 1507
rect 3046 1503 3049 1507
rect 3054 1503 3056 1507
rect 3030 1302 3033 1328
rect 3040 1303 3042 1307
rect 3046 1303 3049 1307
rect 3054 1303 3056 1307
rect 3062 1222 3065 1548
rect 3070 1472 3073 1548
rect 3070 1242 3073 1468
rect 3030 1132 3033 1158
rect 3040 1103 3042 1107
rect 3046 1103 3049 1107
rect 3054 1103 3056 1107
rect 3030 892 3033 1088
rect 3062 1062 3065 1098
rect 3054 932 3057 1018
rect 3066 928 3070 931
rect 3040 903 3042 907
rect 3046 903 3049 907
rect 3054 903 3056 907
rect 3038 888 3046 891
rect 3030 482 3033 848
rect 3038 732 3041 888
rect 3078 742 3081 1548
rect 3086 1332 3089 1378
rect 3086 1262 3089 1308
rect 3110 1272 3113 1338
rect 3126 1212 3129 1508
rect 3134 1372 3137 1618
rect 3158 1572 3161 1588
rect 3142 1492 3145 1528
rect 3134 1252 3137 1348
rect 3142 1292 3145 1488
rect 3086 952 3089 958
rect 3094 952 3097 1168
rect 3106 1138 3110 1141
rect 3040 703 3042 707
rect 3046 703 3049 707
rect 3054 703 3056 707
rect 3066 668 3070 671
rect 3042 638 3046 641
rect 3070 592 3073 658
rect 3040 503 3042 507
rect 3046 503 3049 507
rect 3054 503 3056 507
rect 2930 68 2934 71
rect 2854 52 2857 68
rect 2950 41 2953 88
rect 2966 52 2969 158
rect 2974 72 2977 78
rect 2982 52 2985 198
rect 2950 38 2958 41
rect 2966 32 2969 38
rect 2974 32 2977 38
rect 2990 22 2993 218
rect 3014 112 3017 148
rect 3022 112 3025 138
rect 3030 102 3033 458
rect 3070 422 3073 438
rect 3038 352 3041 368
rect 3078 362 3081 738
rect 3086 512 3089 878
rect 3094 812 3097 948
rect 3102 912 3105 1008
rect 3094 742 3097 758
rect 3102 682 3105 848
rect 3118 842 3121 848
rect 3166 842 3169 1608
rect 3174 1532 3177 1618
rect 3174 842 3177 1528
rect 3182 1202 3185 1518
rect 3190 1362 3193 1788
rect 3198 1612 3201 1748
rect 3214 1692 3217 1708
rect 3210 1688 3214 1691
rect 3210 1458 3214 1461
rect 3214 1282 3217 1448
rect 3182 1152 3185 1158
rect 3182 1072 3185 1118
rect 3166 762 3169 778
rect 3154 688 3158 691
rect 3094 482 3097 558
rect 3102 502 3105 578
rect 3162 548 3166 551
rect 3178 548 3182 551
rect 3078 352 3081 358
rect 3102 342 3105 498
rect 3110 468 3118 471
rect 3110 452 3113 468
rect 3134 462 3137 468
rect 3142 462 3145 528
rect 3182 452 3185 498
rect 3158 372 3161 388
rect 3130 348 3134 351
rect 3138 338 3142 341
rect 3118 332 3121 338
rect 3182 322 3185 428
rect 3042 318 3046 321
rect 3040 303 3042 307
rect 3046 303 3049 307
rect 3054 303 3056 307
rect 3050 188 3054 191
rect 3040 103 3042 107
rect 3046 103 3049 107
rect 3054 103 3056 107
rect 3038 72 3041 78
rect 3030 52 3033 68
rect 3070 62 3073 128
rect 3078 12 3081 268
rect 3190 212 3193 1278
rect 3214 1042 3217 1098
rect 3222 1082 3225 1928
rect 3230 1502 3233 1888
rect 3254 1692 3257 1868
rect 3250 1458 3254 1461
rect 3270 1392 3273 1928
rect 3278 1922 3281 1958
rect 3278 1392 3281 1668
rect 3294 1642 3297 2118
rect 3302 1792 3305 2068
rect 3334 1962 3337 2348
rect 3342 2222 3345 2468
rect 3350 2452 3353 2848
rect 3350 2342 3353 2358
rect 3342 2152 3345 2158
rect 3346 2128 3350 2131
rect 3358 2072 3361 3198
rect 3366 3012 3369 3258
rect 3366 2862 3369 2868
rect 3366 2402 3369 2478
rect 3366 2342 3369 2358
rect 3366 2222 3369 2288
rect 3354 2048 3358 2051
rect 3326 1822 3329 1828
rect 3330 1648 3334 1651
rect 3310 1642 3313 1648
rect 3230 1342 3233 1378
rect 3274 1338 3278 1341
rect 3210 948 3214 951
rect 3222 932 3225 1078
rect 3230 942 3233 948
rect 3238 942 3241 978
rect 3226 848 3230 851
rect 3222 702 3225 728
rect 3206 642 3209 688
rect 3214 672 3217 688
rect 3198 612 3201 638
rect 3198 492 3201 608
rect 3222 482 3225 678
rect 3246 662 3249 668
rect 3234 548 3238 551
rect 3202 348 3206 351
rect 3230 342 3233 538
rect 3242 388 3249 391
rect 3246 292 3249 388
rect 3254 212 3257 1198
rect 3278 1122 3281 1248
rect 3278 1082 3281 1088
rect 3274 938 3278 941
rect 3262 322 3265 328
rect 3094 102 3097 188
rect 3102 122 3105 148
rect 3110 142 3113 148
rect 3182 132 3185 148
rect 3102 92 3105 98
rect 3134 51 3137 118
rect 3134 48 3142 51
rect 3254 42 3257 208
rect 3286 81 3289 1418
rect 3294 742 3297 1478
rect 3302 1292 3305 1328
rect 3310 1322 3313 1358
rect 3318 1292 3321 1458
rect 3302 1132 3305 1138
rect 3294 652 3297 738
rect 3294 552 3297 648
rect 3302 122 3305 1118
rect 3310 1112 3313 1168
rect 3326 1122 3329 1598
rect 3342 1532 3345 1958
rect 3350 1682 3353 1798
rect 3358 1672 3361 1688
rect 3366 1482 3369 1688
rect 3374 1472 3377 3258
rect 3382 2622 3385 2738
rect 3382 2312 3385 2338
rect 3382 1522 3385 2298
rect 3390 1792 3393 3268
rect 3390 1652 3393 1658
rect 3334 1362 3337 1468
rect 3334 1332 3337 1338
rect 3342 1272 3345 1458
rect 3350 1438 3358 1441
rect 3350 1322 3353 1438
rect 3358 1342 3361 1418
rect 3390 1402 3393 1558
rect 3362 1328 3366 1331
rect 3350 1062 3353 1318
rect 3358 1132 3361 1308
rect 3374 1142 3377 1148
rect 3310 132 3313 1058
rect 3346 1048 3350 1051
rect 3346 968 3350 971
rect 3358 492 3361 1128
rect 3382 1062 3385 1128
rect 3370 1048 3374 1051
rect 3330 468 3334 471
rect 3318 152 3321 468
rect 3326 392 3329 448
rect 3318 132 3321 148
rect 3286 78 3294 81
rect 3310 72 3313 118
rect 3326 102 3329 378
rect 3322 68 3326 71
rect 3334 12 3337 278
rect 3342 142 3345 458
rect 3350 132 3353 138
rect 3358 132 3361 488
rect 3366 182 3369 1028
rect 3374 642 3377 968
rect 3382 952 3385 1058
rect 3390 642 3393 1388
rect 3390 182 3393 188
rect 3398 162 3401 3258
rect 3422 2602 3425 2938
rect 3406 2352 3409 2358
rect 3414 1992 3417 2588
rect 3422 2292 3425 2458
rect 3406 1742 3409 1768
rect 3414 1742 3417 1988
rect 3430 1782 3433 2348
rect 3406 1552 3409 1678
rect 3406 1362 3409 1468
rect 3406 1332 3409 1338
rect 3414 1292 3417 1728
rect 3422 1662 3425 1768
rect 3438 1752 3441 3268
rect 3458 3258 3462 3261
rect 3450 3248 3454 3251
rect 3446 2742 3449 2888
rect 3446 2342 3449 2738
rect 3454 2352 3457 2788
rect 3458 2338 3462 2341
rect 3446 2112 3449 2148
rect 3454 2082 3457 2168
rect 3422 1482 3425 1568
rect 3422 1332 3425 1448
rect 3430 1412 3433 1518
rect 3430 1322 3433 1338
rect 3426 1258 3433 1261
rect 3430 1042 3433 1258
rect 3422 952 3425 958
rect 3410 478 3414 481
rect 3438 472 3441 1748
rect 3462 1582 3465 2328
rect 3470 1702 3473 3138
rect 3478 2362 3481 2778
rect 3486 2172 3489 2878
rect 3486 2102 3489 2138
rect 3494 2091 3497 3138
rect 3486 2088 3497 2091
rect 3470 1642 3473 1648
rect 3446 1512 3449 1548
rect 3454 592 3457 1348
rect 3462 1302 3465 1508
rect 3470 1032 3473 1538
rect 3478 1342 3481 1718
rect 3478 1282 3481 1328
rect 3486 1272 3489 2088
rect 3502 1912 3505 3228
rect 3494 1112 3497 1738
rect 3502 1732 3505 1898
rect 3502 1332 3505 1728
rect 3510 1662 3513 2978
rect 3518 1702 3521 2898
rect 3526 2592 3529 2868
rect 3534 2442 3537 2898
rect 3542 2752 3545 2958
rect 3526 1712 3529 1898
rect 3534 1742 3537 1908
rect 3542 1842 3545 1868
rect 3510 1482 3513 1578
rect 3510 982 3513 998
rect 3466 958 3470 961
rect 3406 342 3409 408
rect 3430 362 3433 398
rect 3422 322 3425 328
rect 3430 262 3433 358
rect 3366 132 3369 138
rect 3342 82 3345 98
rect 3346 68 3350 71
rect 3398 52 3401 158
rect 3438 82 3441 468
rect 3454 112 3457 588
rect 3462 82 3465 778
rect 3474 348 3478 351
rect 3518 142 3521 1678
rect 3526 1482 3529 1688
rect 3534 1562 3537 1738
rect 3550 1722 3553 3248
rect 3558 2062 3561 2068
rect 3558 1772 3561 1778
rect 3558 1752 3561 1758
rect 3558 1672 3561 1678
rect 3526 1462 3529 1468
rect 3526 992 3529 998
rect 3534 772 3537 1548
rect 3542 972 3545 1658
rect 3558 1552 3561 1588
rect 3526 122 3529 508
rect 3482 68 3486 71
rect 3550 62 3553 1548
rect 3558 1142 3561 1148
rect 2414 8 2422 11
rect 480 3 482 7
rect 486 3 489 7
rect 494 3 496 7
rect 1512 3 1514 7
rect 1518 3 1521 7
rect 1526 3 1528 7
rect 2536 3 2538 7
rect 2542 3 2545 7
rect 2550 3 2552 7
<< m5contact >>
rect 994 3303 998 3307
rect 1001 3303 1002 3307
rect 1002 3303 1005 3307
rect 2026 3303 2030 3307
rect 2033 3303 2034 3307
rect 2034 3303 2037 3307
rect 3042 3303 3046 3307
rect 3049 3303 3050 3307
rect 3050 3303 3053 3307
rect 1142 3298 1146 3302
rect 482 3203 486 3207
rect 489 3203 490 3207
rect 490 3203 493 3207
rect 166 3058 170 3062
rect 6 2558 10 2562
rect 22 2368 26 2372
rect 6 2358 10 2362
rect 6 2338 10 2342
rect 182 2748 186 2752
rect 14 2238 18 2242
rect 102 2448 106 2452
rect 198 2528 202 2532
rect 182 2518 186 2522
rect 78 1978 82 1982
rect 6 978 10 982
rect 118 858 122 862
rect 134 1738 138 1742
rect 134 1488 138 1492
rect 230 2918 234 2922
rect 238 2868 242 2872
rect 286 2878 290 2882
rect 294 2858 298 2862
rect 614 3258 618 3262
rect 342 3058 346 3062
rect 574 3058 578 3062
rect 334 3038 338 3042
rect 438 3038 442 3042
rect 374 2858 378 2862
rect 278 2848 282 2852
rect 350 2848 354 2852
rect 390 2878 394 2882
rect 382 2788 386 2792
rect 326 2748 330 2752
rect 278 2548 282 2552
rect 214 2488 218 2492
rect 206 2178 210 2182
rect 230 2148 234 2152
rect 174 2128 178 2132
rect 166 1858 170 1862
rect 166 1738 170 1742
rect 158 1518 162 1522
rect 190 1888 194 1892
rect 174 838 178 842
rect 126 658 130 662
rect 390 2638 394 2642
rect 374 2518 378 2522
rect 286 2378 290 2382
rect 270 2078 274 2082
rect 230 1788 234 1792
rect 238 1748 242 1752
rect 302 2038 306 2042
rect 270 1828 274 1832
rect 342 2278 346 2282
rect 286 1748 290 1752
rect 278 1678 282 1682
rect 214 1358 218 1362
rect 230 1358 234 1362
rect 206 1248 210 1252
rect 198 618 202 622
rect 110 268 114 272
rect 198 168 202 172
rect 246 1248 250 1252
rect 230 1228 234 1232
rect 230 1058 234 1062
rect 246 708 250 712
rect 238 538 242 542
rect 246 508 250 512
rect 126 138 130 142
rect 318 1708 322 1712
rect 310 1688 314 1692
rect 286 1528 290 1532
rect 366 2318 370 2322
rect 366 2228 370 2232
rect 334 1698 338 1702
rect 334 1578 338 1582
rect 334 1428 338 1432
rect 482 3003 486 3007
rect 489 3003 490 3007
rect 490 3003 493 3007
rect 446 2718 450 2722
rect 510 2868 514 2872
rect 482 2803 486 2807
rect 489 2803 490 2807
rect 490 2803 493 2807
rect 438 2588 442 2592
rect 438 2518 442 2522
rect 502 2708 506 2712
rect 518 2658 522 2662
rect 478 2638 482 2642
rect 482 2603 486 2607
rect 489 2603 490 2607
rect 490 2603 493 2607
rect 470 2578 474 2582
rect 462 2548 466 2552
rect 550 2878 554 2882
rect 566 2768 570 2772
rect 534 2728 538 2732
rect 526 2538 530 2542
rect 534 2528 538 2532
rect 614 3058 618 3062
rect 470 2478 474 2482
rect 582 2558 586 2562
rect 614 2588 618 2592
rect 614 2548 618 2552
rect 614 2508 618 2512
rect 598 2448 602 2452
rect 414 2428 418 2432
rect 502 2428 506 2432
rect 582 2428 586 2432
rect 502 2408 506 2412
rect 390 2348 394 2352
rect 406 2318 410 2322
rect 406 1978 410 1982
rect 454 2338 458 2342
rect 482 2403 486 2407
rect 489 2403 490 2407
rect 490 2403 493 2407
rect 526 2388 530 2392
rect 718 3048 722 3052
rect 750 2938 754 2942
rect 814 2948 818 2952
rect 838 2928 842 2932
rect 846 2918 850 2922
rect 774 2878 778 2882
rect 982 3138 986 3142
rect 902 3118 906 3122
rect 994 3103 998 3107
rect 1001 3103 1002 3107
rect 1002 3103 1005 3107
rect 910 3088 914 3092
rect 942 3078 946 3082
rect 918 2938 922 2942
rect 862 2918 866 2922
rect 910 2868 914 2872
rect 654 2718 658 2722
rect 646 2668 650 2672
rect 646 2648 650 2652
rect 694 2738 698 2742
rect 742 2718 746 2722
rect 750 2708 754 2712
rect 774 2658 778 2662
rect 718 2648 722 2652
rect 774 2558 778 2562
rect 654 2458 658 2462
rect 654 2438 658 2442
rect 574 2368 578 2372
rect 542 2328 546 2332
rect 558 2348 562 2352
rect 574 2338 578 2342
rect 518 2208 522 2212
rect 482 2203 486 2207
rect 489 2203 490 2207
rect 490 2203 493 2207
rect 566 2258 570 2262
rect 622 2358 626 2362
rect 670 2418 674 2422
rect 590 2318 594 2322
rect 606 2318 610 2322
rect 590 2248 594 2252
rect 574 2238 578 2242
rect 582 2168 586 2172
rect 550 2158 554 2162
rect 582 2148 586 2152
rect 598 2148 602 2152
rect 526 2078 530 2082
rect 526 2068 530 2072
rect 470 2028 474 2032
rect 482 2003 486 2007
rect 489 2003 490 2007
rect 490 2003 493 2007
rect 470 1978 474 1982
rect 398 1858 402 1862
rect 382 1818 386 1822
rect 366 1718 370 1722
rect 398 1658 402 1662
rect 358 1508 362 1512
rect 350 1478 354 1482
rect 350 1378 354 1382
rect 366 1328 370 1332
rect 302 1248 306 1252
rect 286 838 290 842
rect 278 728 282 732
rect 270 668 274 672
rect 286 528 290 532
rect 278 268 282 272
rect 310 758 314 762
rect 342 858 346 862
rect 350 818 354 822
rect 310 698 314 702
rect 334 688 338 692
rect 302 648 306 652
rect 398 1438 402 1442
rect 534 1978 538 1982
rect 518 1878 522 1882
rect 558 1868 562 1872
rect 454 1848 458 1852
rect 430 1778 434 1782
rect 482 1803 486 1807
rect 489 1803 490 1807
rect 490 1803 493 1807
rect 454 1768 458 1772
rect 414 1578 418 1582
rect 422 1478 426 1482
rect 414 1308 418 1312
rect 398 1248 402 1252
rect 390 1178 394 1182
rect 398 1148 402 1152
rect 398 968 402 972
rect 390 958 394 962
rect 358 718 362 722
rect 382 638 386 642
rect 366 448 370 452
rect 494 1758 498 1762
rect 494 1648 498 1652
rect 482 1603 486 1607
rect 489 1603 490 1607
rect 490 1603 493 1607
rect 470 1588 474 1592
rect 470 1558 474 1562
rect 446 1478 450 1482
rect 446 1388 450 1392
rect 454 1248 458 1252
rect 446 1238 450 1242
rect 462 1218 466 1222
rect 462 1158 466 1162
rect 438 1048 442 1052
rect 518 1738 522 1742
rect 510 1728 514 1732
rect 482 1403 486 1407
rect 489 1403 490 1407
rect 490 1403 493 1407
rect 482 1203 486 1207
rect 489 1203 490 1207
rect 490 1203 493 1207
rect 542 1708 546 1712
rect 542 1548 546 1552
rect 534 1518 538 1522
rect 518 1358 522 1362
rect 526 1338 530 1342
rect 510 1148 514 1152
rect 502 1038 506 1042
rect 482 1003 486 1007
rect 489 1003 490 1007
rect 490 1003 493 1007
rect 502 978 506 982
rect 470 958 474 962
rect 462 928 466 932
rect 462 848 466 852
rect 454 768 458 772
rect 422 618 426 622
rect 398 548 402 552
rect 406 488 410 492
rect 454 638 458 642
rect 438 518 442 522
rect 454 478 458 482
rect 482 803 486 807
rect 489 803 490 807
rect 490 803 493 807
rect 482 603 486 607
rect 489 603 490 607
rect 490 603 493 607
rect 550 1538 554 1542
rect 542 788 546 792
rect 542 738 546 742
rect 510 588 514 592
rect 502 558 506 562
rect 470 538 474 542
rect 598 2068 602 2072
rect 598 2058 602 2062
rect 590 1858 594 1862
rect 590 1808 594 1812
rect 574 1788 578 1792
rect 566 1548 570 1552
rect 590 1718 594 1722
rect 590 1568 594 1572
rect 574 1528 578 1532
rect 590 1358 594 1362
rect 574 1168 578 1172
rect 558 848 562 852
rect 582 1048 586 1052
rect 574 888 578 892
rect 590 828 594 832
rect 550 548 554 552
rect 518 498 522 502
rect 482 403 486 407
rect 489 403 490 407
rect 490 403 493 407
rect 478 378 482 382
rect 470 328 474 332
rect 390 318 394 322
rect 454 318 458 322
rect 482 203 486 207
rect 489 203 490 207
rect 490 203 493 207
rect 374 108 378 112
rect 366 98 370 102
rect 438 118 442 122
rect 446 108 450 112
rect 350 88 354 92
rect 110 78 114 82
rect 542 328 546 332
rect 566 618 570 622
rect 606 2018 610 2022
rect 614 1938 618 1942
rect 622 1938 626 1942
rect 646 2108 650 2112
rect 662 2328 666 2332
rect 670 2238 674 2242
rect 678 2198 682 2202
rect 726 2408 730 2412
rect 734 2358 738 2362
rect 694 2228 698 2232
rect 686 2188 690 2192
rect 734 2338 738 2342
rect 726 2308 730 2312
rect 710 2278 714 2282
rect 726 2278 730 2282
rect 758 2348 762 2352
rect 726 2188 730 2192
rect 686 2078 690 2082
rect 718 2068 722 2072
rect 654 1998 658 2002
rect 686 1988 690 1992
rect 622 1868 626 1872
rect 654 1828 658 1832
rect 638 1798 642 1802
rect 726 1858 730 1862
rect 694 1828 698 1832
rect 686 1778 690 1782
rect 646 1748 650 1752
rect 694 1748 698 1752
rect 646 1738 650 1742
rect 654 1728 658 1732
rect 622 1668 626 1672
rect 614 1658 618 1662
rect 606 1558 610 1562
rect 630 1598 634 1602
rect 606 1528 610 1532
rect 662 1608 666 1612
rect 630 1458 634 1462
rect 654 1448 658 1452
rect 646 1348 650 1352
rect 614 1278 618 1282
rect 622 1268 626 1272
rect 622 1088 626 1092
rect 614 1068 618 1072
rect 606 988 610 992
rect 622 1048 626 1052
rect 622 938 626 942
rect 678 1678 682 1682
rect 678 1638 682 1642
rect 670 1308 674 1312
rect 654 1258 658 1262
rect 710 1718 714 1722
rect 710 1698 714 1702
rect 726 1738 730 1742
rect 726 1628 730 1632
rect 702 1538 706 1542
rect 694 1478 698 1482
rect 686 1248 690 1252
rect 686 1158 690 1162
rect 670 1138 674 1142
rect 662 1108 666 1112
rect 654 1048 658 1052
rect 654 948 658 952
rect 638 888 642 892
rect 606 758 610 762
rect 606 718 610 722
rect 598 678 602 682
rect 590 658 594 662
rect 598 648 602 652
rect 606 628 610 632
rect 622 818 626 822
rect 670 1028 674 1032
rect 662 808 666 812
rect 654 788 658 792
rect 638 708 642 712
rect 606 438 610 442
rect 590 368 594 372
rect 590 358 594 362
rect 582 338 586 342
rect 590 338 594 342
rect 558 158 562 162
rect 542 148 546 152
rect 566 98 570 102
rect 430 68 434 72
rect 558 58 562 62
rect 486 48 490 52
rect 630 468 634 472
rect 622 418 626 422
rect 614 398 618 402
rect 726 1318 730 1322
rect 726 1208 730 1212
rect 750 2218 754 2222
rect 886 2768 890 2772
rect 870 2758 874 2762
rect 846 2638 850 2642
rect 846 2628 850 2632
rect 838 2568 842 2572
rect 798 2428 802 2432
rect 782 2328 786 2332
rect 774 2168 778 2172
rect 774 2128 778 2132
rect 798 2308 802 2312
rect 830 2458 834 2462
rect 846 2418 850 2422
rect 822 2408 826 2412
rect 750 1528 754 1532
rect 742 1398 746 1402
rect 742 1268 746 1272
rect 750 1198 754 1202
rect 710 1148 714 1152
rect 726 1118 730 1122
rect 710 1098 714 1102
rect 718 1038 722 1042
rect 734 1038 738 1042
rect 742 1028 746 1032
rect 710 918 714 922
rect 718 878 722 882
rect 678 688 682 692
rect 710 838 714 842
rect 670 598 674 602
rect 686 478 690 482
rect 654 358 658 362
rect 622 328 626 332
rect 662 328 666 332
rect 606 238 610 242
rect 630 258 634 262
rect 622 208 626 212
rect 686 228 690 232
rect 662 148 666 152
rect 670 108 674 112
rect 622 98 626 102
rect 694 218 698 222
rect 694 188 698 192
rect 742 898 746 902
rect 734 778 738 782
rect 718 708 722 712
rect 718 698 722 702
rect 710 688 714 692
rect 718 648 722 652
rect 798 2058 802 2062
rect 790 1778 794 1782
rect 766 1688 770 1692
rect 782 1678 786 1682
rect 774 1628 778 1632
rect 774 1618 778 1622
rect 782 1578 786 1582
rect 782 1558 786 1562
rect 782 1278 786 1282
rect 782 1078 786 1082
rect 798 1248 802 1252
rect 798 1008 802 1012
rect 782 918 786 922
rect 758 848 762 852
rect 742 558 746 562
rect 734 548 738 552
rect 710 478 714 482
rect 750 388 754 392
rect 702 178 706 182
rect 718 178 722 182
rect 766 788 770 792
rect 766 708 770 712
rect 798 888 802 892
rect 798 868 802 872
rect 814 2148 818 2152
rect 814 1738 818 1742
rect 870 2648 874 2652
rect 878 2588 882 2592
rect 990 2938 994 2942
rect 998 2928 1002 2932
rect 1014 2928 1018 2932
rect 974 2918 978 2922
rect 994 2903 998 2907
rect 1001 2903 1002 2907
rect 1002 2903 1005 2907
rect 934 2888 938 2892
rect 950 2758 954 2762
rect 910 2658 914 2662
rect 878 2468 882 2472
rect 886 2418 890 2422
rect 854 2248 858 2252
rect 854 2188 858 2192
rect 902 2368 906 2372
rect 902 2358 906 2362
rect 942 2658 946 2662
rect 942 2638 946 2642
rect 926 2588 930 2592
rect 950 2538 954 2542
rect 942 2508 946 2512
rect 934 2488 938 2492
rect 886 2338 890 2342
rect 878 2038 882 2042
rect 846 2008 850 2012
rect 870 1728 874 1732
rect 854 1718 858 1722
rect 862 1668 866 1672
rect 862 1518 866 1522
rect 870 1408 874 1412
rect 854 1368 858 1372
rect 830 1328 834 1332
rect 854 1308 858 1312
rect 854 1288 858 1292
rect 870 1278 874 1282
rect 862 1268 866 1272
rect 846 1258 850 1262
rect 846 1228 850 1232
rect 870 1218 874 1222
rect 830 1178 834 1182
rect 846 1168 850 1172
rect 822 1148 826 1152
rect 838 1148 842 1152
rect 838 1128 842 1132
rect 814 1098 818 1102
rect 822 968 826 972
rect 782 798 786 802
rect 790 748 794 752
rect 782 638 786 642
rect 790 588 794 592
rect 798 578 802 582
rect 766 488 770 492
rect 774 488 778 492
rect 774 378 778 382
rect 742 168 746 172
rect 774 168 778 172
rect 726 138 730 142
rect 766 138 770 142
rect 734 128 738 132
rect 686 88 690 92
rect 702 88 706 92
rect 798 308 802 312
rect 758 78 762 82
rect 782 78 786 82
rect 814 808 818 812
rect 838 1048 842 1052
rect 846 1048 850 1052
rect 870 1128 874 1132
rect 870 1088 874 1092
rect 846 998 850 1002
rect 838 958 842 962
rect 862 968 866 972
rect 870 968 874 972
rect 838 848 842 852
rect 814 558 818 562
rect 830 738 834 742
rect 838 738 842 742
rect 830 658 834 662
rect 838 548 842 552
rect 822 538 826 542
rect 862 908 866 912
rect 870 868 874 872
rect 886 1568 890 1572
rect 886 1518 890 1522
rect 886 1478 890 1482
rect 862 838 866 842
rect 878 728 882 732
rect 878 718 882 722
rect 886 698 890 702
rect 886 648 890 652
rect 854 528 858 532
rect 878 518 882 522
rect 846 408 850 412
rect 846 308 850 312
rect 806 248 810 252
rect 886 428 890 432
rect 886 218 890 222
rect 878 188 882 192
rect 838 168 842 172
rect 830 158 834 162
rect 846 158 850 162
rect 710 48 714 52
rect 702 38 706 42
rect 790 38 794 42
rect 726 28 730 32
rect 646 18 650 22
rect 814 98 818 102
rect 838 78 842 82
rect 910 1398 914 1402
rect 910 1148 914 1152
rect 910 1068 914 1072
rect 910 1018 914 1022
rect 910 998 914 1002
rect 910 668 914 672
rect 910 658 914 662
rect 910 578 914 582
rect 910 358 914 362
rect 926 2148 930 2152
rect 926 2108 930 2112
rect 934 2088 938 2092
rect 994 2703 998 2707
rect 1001 2703 1002 2707
rect 1002 2703 1005 2707
rect 998 2688 1002 2692
rect 974 2568 978 2572
rect 1006 2518 1010 2522
rect 994 2503 998 2507
rect 1001 2503 1002 2507
rect 1002 2503 1005 2507
rect 974 2488 978 2492
rect 966 2388 970 2392
rect 958 2348 962 2352
rect 950 2188 954 2192
rect 1054 3238 1058 3242
rect 1062 2938 1066 2942
rect 1102 3188 1106 3192
rect 1118 3118 1122 3122
rect 1118 3078 1122 3082
rect 1046 2728 1050 2732
rect 1054 2648 1058 2652
rect 1030 2538 1034 2542
rect 1022 2388 1026 2392
rect 1006 2348 1010 2352
rect 994 2303 998 2307
rect 1001 2303 1002 2307
rect 1002 2303 1005 2307
rect 982 2288 986 2292
rect 1014 2278 1018 2282
rect 990 2158 994 2162
rect 974 2138 978 2142
rect 998 2128 1002 2132
rect 966 2048 970 2052
rect 942 1948 946 1952
rect 934 1898 938 1902
rect 934 1718 938 1722
rect 926 1708 930 1712
rect 950 1928 954 1932
rect 926 1208 930 1212
rect 966 1968 970 1972
rect 950 1598 954 1602
rect 942 1558 946 1562
rect 994 2103 998 2107
rect 1001 2103 1002 2107
rect 1002 2103 1005 2107
rect 974 1938 978 1942
rect 994 1903 998 1907
rect 1001 1903 1002 1907
rect 1002 1903 1005 1907
rect 998 1878 1002 1882
rect 966 1698 970 1702
rect 990 1768 994 1772
rect 994 1703 998 1707
rect 1001 1703 1002 1707
rect 1002 1703 1005 1707
rect 974 1658 978 1662
rect 966 1648 970 1652
rect 958 1538 962 1542
rect 942 1518 946 1522
rect 1006 1598 1010 1602
rect 994 1503 998 1507
rect 1001 1503 1002 1507
rect 1002 1503 1005 1507
rect 982 1478 986 1482
rect 998 1458 1002 1462
rect 982 1448 986 1452
rect 982 1398 986 1402
rect 950 1368 954 1372
rect 966 1348 970 1352
rect 982 1348 986 1352
rect 966 1338 970 1342
rect 942 1328 946 1332
rect 942 1268 946 1272
rect 974 1328 978 1332
rect 966 1318 970 1322
rect 974 1308 978 1312
rect 1006 1448 1010 1452
rect 998 1418 1002 1422
rect 998 1408 1002 1412
rect 1006 1408 1010 1412
rect 990 1318 994 1322
rect 1006 1318 1010 1322
rect 994 1303 998 1307
rect 1001 1303 1002 1307
rect 1002 1303 1005 1307
rect 950 1258 954 1262
rect 966 1258 970 1262
rect 998 1248 1002 1252
rect 942 1208 946 1212
rect 990 1208 994 1212
rect 950 1168 954 1172
rect 974 1188 978 1192
rect 926 1138 930 1142
rect 926 848 930 852
rect 982 1108 986 1112
rect 994 1103 998 1107
rect 1001 1103 1002 1107
rect 1002 1103 1005 1107
rect 966 1088 970 1092
rect 958 978 962 982
rect 982 1048 986 1052
rect 974 1018 978 1022
rect 1006 1018 1010 1022
rect 982 958 986 962
rect 974 938 978 942
rect 982 908 986 912
rect 994 903 998 907
rect 1001 903 1002 907
rect 1002 903 1005 907
rect 942 868 946 872
rect 966 868 970 872
rect 958 858 962 862
rect 998 868 1002 872
rect 966 778 970 782
rect 990 758 994 762
rect 934 638 938 642
rect 926 598 930 602
rect 934 578 938 582
rect 934 548 938 552
rect 974 708 978 712
rect 950 678 954 682
rect 942 508 946 512
rect 950 448 954 452
rect 994 703 998 707
rect 1001 703 1002 707
rect 1002 703 1005 707
rect 982 678 986 682
rect 974 638 978 642
rect 966 558 970 562
rect 1006 578 1010 582
rect 994 503 998 507
rect 1001 503 1002 507
rect 1002 503 1005 507
rect 1006 438 1010 442
rect 934 358 938 362
rect 958 358 962 362
rect 926 278 930 282
rect 926 228 930 232
rect 934 208 938 212
rect 950 178 954 182
rect 926 168 930 172
rect 870 68 874 72
rect 942 118 946 122
rect 926 78 930 82
rect 994 303 998 307
rect 1001 303 1002 307
rect 1002 303 1005 307
rect 1054 2528 1058 2532
rect 1070 2848 1074 2852
rect 1038 2498 1042 2502
rect 1062 2488 1066 2492
rect 1038 2448 1042 2452
rect 1030 2338 1034 2342
rect 1022 2018 1026 2022
rect 1022 1708 1026 1712
rect 1086 2568 1090 2572
rect 1078 2558 1082 2562
rect 1062 2268 1066 2272
rect 1070 2198 1074 2202
rect 1038 2018 1042 2022
rect 1046 1918 1050 1922
rect 1126 2908 1130 2912
rect 1118 2878 1122 2882
rect 1150 2988 1154 2992
rect 1182 2948 1186 2952
rect 1134 2868 1138 2872
rect 1126 2668 1130 2672
rect 1190 2748 1194 2752
rect 1158 2658 1162 2662
rect 1150 2628 1154 2632
rect 1334 3138 1338 3142
rect 1342 3088 1346 3092
rect 1326 2928 1330 2932
rect 1294 2888 1298 2892
rect 1238 2848 1242 2852
rect 1222 2748 1226 2752
rect 1222 2698 1226 2702
rect 1214 2678 1218 2682
rect 1206 2658 1210 2662
rect 1134 2568 1138 2572
rect 1150 2568 1154 2572
rect 1118 2548 1122 2552
rect 1126 2548 1130 2552
rect 1102 2488 1106 2492
rect 1102 2468 1106 2472
rect 1118 2438 1122 2442
rect 1086 2338 1090 2342
rect 1118 2298 1122 2302
rect 1086 2078 1090 2082
rect 1102 2218 1106 2222
rect 1102 2068 1106 2072
rect 1102 2018 1106 2022
rect 1086 1928 1090 1932
rect 1094 1868 1098 1872
rect 1078 1828 1082 1832
rect 1062 1768 1066 1772
rect 1070 1768 1074 1772
rect 1054 1728 1058 1732
rect 1038 1708 1042 1712
rect 1046 1708 1050 1712
rect 1038 1668 1042 1672
rect 1062 1668 1066 1672
rect 1054 1658 1058 1662
rect 1054 1578 1058 1582
rect 1054 1548 1058 1552
rect 1030 1538 1034 1542
rect 1030 1468 1034 1472
rect 1062 1508 1066 1512
rect 1022 1458 1026 1462
rect 1030 1458 1034 1462
rect 1062 1448 1066 1452
rect 1046 1418 1050 1422
rect 1054 1418 1058 1422
rect 1030 1408 1034 1412
rect 1022 1348 1026 1352
rect 1030 1338 1034 1342
rect 1046 1348 1050 1352
rect 1038 1308 1042 1312
rect 1030 1268 1034 1272
rect 1022 1248 1026 1252
rect 1022 1208 1026 1212
rect 1022 1158 1026 1162
rect 1038 1248 1042 1252
rect 1062 1378 1066 1382
rect 1086 1788 1090 1792
rect 1094 1778 1098 1782
rect 1134 2448 1138 2452
rect 1158 2378 1162 2382
rect 1150 2368 1154 2372
rect 1126 2238 1130 2242
rect 1190 2328 1194 2332
rect 1174 2258 1178 2262
rect 1182 2228 1186 2232
rect 1214 2558 1218 2562
rect 1222 2508 1226 2512
rect 1326 2718 1330 2722
rect 1318 2708 1322 2712
rect 1326 2678 1330 2682
rect 1302 2638 1306 2642
rect 1254 2548 1258 2552
rect 1278 2538 1282 2542
rect 1238 2458 1242 2462
rect 1230 2368 1234 2372
rect 1214 2318 1218 2322
rect 1262 2478 1266 2482
rect 1294 2438 1298 2442
rect 1270 2388 1274 2392
rect 1270 2378 1274 2382
rect 1278 2368 1282 2372
rect 1246 2308 1250 2312
rect 1294 2308 1298 2312
rect 1254 2268 1258 2272
rect 1238 2188 1242 2192
rect 1230 2118 1234 2122
rect 1118 1828 1122 1832
rect 1142 1858 1146 1862
rect 1142 1778 1146 1782
rect 1134 1728 1138 1732
rect 1118 1668 1122 1672
rect 1134 1648 1138 1652
rect 1134 1618 1138 1622
rect 1134 1598 1138 1602
rect 1102 1578 1106 1582
rect 1126 1578 1130 1582
rect 1094 1418 1098 1422
rect 1086 1368 1090 1372
rect 1094 1368 1098 1372
rect 1070 1318 1074 1322
rect 1046 1178 1050 1182
rect 1118 1488 1122 1492
rect 1158 1868 1162 1872
rect 1158 1728 1162 1732
rect 1182 1898 1186 1902
rect 1286 2288 1290 2292
rect 1206 1878 1210 1882
rect 1158 1708 1162 1712
rect 1166 1668 1170 1672
rect 1198 1718 1202 1722
rect 1206 1718 1210 1722
rect 1190 1678 1194 1682
rect 1166 1658 1170 1662
rect 1142 1548 1146 1552
rect 1174 1598 1178 1602
rect 1166 1558 1170 1562
rect 1158 1518 1162 1522
rect 1198 1588 1202 1592
rect 1254 1948 1258 1952
rect 1270 1888 1274 1892
rect 1310 2088 1314 2092
rect 1310 2018 1314 2022
rect 1254 1788 1258 1792
rect 1246 1768 1250 1772
rect 1238 1738 1242 1742
rect 1238 1708 1242 1712
rect 1182 1488 1186 1492
rect 1142 1468 1146 1472
rect 1134 1448 1138 1452
rect 1118 1318 1122 1322
rect 1110 1278 1114 1282
rect 1086 1258 1090 1262
rect 1094 1248 1098 1252
rect 1102 1238 1106 1242
rect 1110 1238 1114 1242
rect 1150 1398 1154 1402
rect 1158 1398 1162 1402
rect 1158 1318 1162 1322
rect 1150 1308 1154 1312
rect 1118 1188 1122 1192
rect 1094 1168 1098 1172
rect 1118 1168 1122 1172
rect 1062 1158 1066 1162
rect 1070 1148 1074 1152
rect 1030 1108 1034 1112
rect 1030 1078 1034 1082
rect 1038 1078 1042 1082
rect 1022 1058 1026 1062
rect 1062 1088 1066 1092
rect 1022 968 1026 972
rect 1086 1138 1090 1142
rect 1070 998 1074 1002
rect 1046 958 1050 962
rect 1054 948 1058 952
rect 1038 898 1042 902
rect 1062 938 1066 942
rect 1046 878 1050 882
rect 1110 1138 1114 1142
rect 1126 1128 1130 1132
rect 1134 1128 1138 1132
rect 1126 1118 1130 1122
rect 1110 1088 1114 1092
rect 1150 1148 1154 1152
rect 1142 1118 1146 1122
rect 1134 1108 1138 1112
rect 1142 1108 1146 1112
rect 1158 1088 1162 1092
rect 1142 1068 1146 1072
rect 1150 1068 1154 1072
rect 1078 938 1082 942
rect 1078 708 1082 712
rect 1070 698 1074 702
rect 1022 658 1026 662
rect 1118 1048 1122 1052
rect 1126 1048 1130 1052
rect 1126 968 1130 972
rect 1110 958 1114 962
rect 1158 1058 1162 1062
rect 1142 908 1146 912
rect 1150 908 1154 912
rect 1190 1458 1194 1462
rect 1230 1538 1234 1542
rect 1262 1598 1266 1602
rect 1262 1588 1266 1592
rect 1254 1578 1258 1582
rect 1262 1528 1266 1532
rect 1278 1688 1282 1692
rect 1366 2768 1370 2772
rect 1534 3268 1538 3272
rect 1422 3258 1426 3262
rect 1406 2818 1410 2822
rect 1422 2738 1426 2742
rect 1358 2698 1362 2702
rect 1398 2698 1402 2702
rect 1422 2698 1426 2702
rect 1398 2588 1402 2592
rect 1358 2498 1362 2502
rect 1366 2428 1370 2432
rect 1350 2408 1354 2412
rect 1350 2318 1354 2322
rect 1406 2538 1410 2542
rect 1406 2458 1410 2462
rect 1390 2418 1394 2422
rect 1382 2098 1386 2102
rect 1366 1958 1370 1962
rect 1374 1848 1378 1852
rect 1326 1838 1330 1842
rect 1334 1828 1338 1832
rect 1342 1828 1346 1832
rect 1310 1768 1314 1772
rect 1310 1758 1314 1762
rect 1294 1738 1298 1742
rect 1294 1678 1298 1682
rect 1294 1658 1298 1662
rect 1294 1598 1298 1602
rect 1294 1578 1298 1582
rect 1286 1558 1290 1562
rect 1278 1498 1282 1502
rect 1286 1498 1290 1502
rect 1206 1458 1210 1462
rect 1230 1448 1234 1452
rect 1198 1418 1202 1422
rect 1214 1368 1218 1372
rect 1230 1368 1234 1372
rect 1206 1338 1210 1342
rect 1206 1268 1210 1272
rect 1206 1238 1210 1242
rect 1190 1188 1194 1192
rect 1174 1118 1178 1122
rect 1190 1098 1194 1102
rect 1174 1008 1178 1012
rect 1182 988 1186 992
rect 1182 938 1186 942
rect 1166 888 1170 892
rect 1118 878 1122 882
rect 1110 858 1114 862
rect 1078 678 1082 682
rect 1038 638 1042 642
rect 1054 638 1058 642
rect 1030 598 1034 602
rect 1046 578 1050 582
rect 1022 508 1026 512
rect 1030 318 1034 322
rect 1022 308 1026 312
rect 1022 258 1026 262
rect 982 168 986 172
rect 1022 108 1026 112
rect 994 103 998 107
rect 1001 103 1002 107
rect 1002 103 1005 107
rect 1006 58 1010 62
rect 1038 48 1042 52
rect 1014 18 1018 22
rect 1086 588 1090 592
rect 1142 828 1146 832
rect 1150 828 1154 832
rect 1166 818 1170 822
rect 1158 788 1162 792
rect 1134 738 1138 742
rect 1158 748 1162 752
rect 1142 698 1146 702
rect 1134 688 1138 692
rect 1126 668 1130 672
rect 1110 608 1114 612
rect 1102 598 1106 602
rect 1110 578 1114 582
rect 1134 578 1138 582
rect 1182 768 1186 772
rect 1182 698 1186 702
rect 1166 688 1170 692
rect 1142 558 1146 562
rect 1102 548 1106 552
rect 1094 518 1098 522
rect 1142 538 1146 542
rect 1110 328 1114 332
rect 1110 278 1114 282
rect 1102 258 1106 262
rect 1182 648 1186 652
rect 1206 1118 1210 1122
rect 1198 1008 1202 1012
rect 1230 1338 1234 1342
rect 1222 1158 1226 1162
rect 1246 1458 1250 1462
rect 1278 1478 1282 1482
rect 1286 1478 1290 1482
rect 1270 1458 1274 1462
rect 1262 1448 1266 1452
rect 1254 1428 1258 1432
rect 1262 1428 1266 1432
rect 1246 1408 1250 1412
rect 1270 1348 1274 1352
rect 1238 1278 1242 1282
rect 1238 1268 1242 1272
rect 1262 1268 1266 1272
rect 1326 1708 1330 1712
rect 1302 1388 1306 1392
rect 1294 1348 1298 1352
rect 1318 1558 1322 1562
rect 1318 1498 1322 1502
rect 1318 1478 1322 1482
rect 1358 1758 1362 1762
rect 1406 2418 1410 2422
rect 1414 2278 1418 2282
rect 1446 3138 1450 3142
rect 1502 3238 1506 3242
rect 1514 3203 1518 3207
rect 1521 3203 1522 3207
rect 1522 3203 1525 3207
rect 1478 3048 1482 3052
rect 1462 3038 1466 3042
rect 1454 3018 1458 3022
rect 1478 2938 1482 2942
rect 1494 3028 1498 3032
rect 1514 3003 1518 3007
rect 1521 3003 1522 3007
rect 1522 3003 1525 3007
rect 1514 2803 1518 2807
rect 1521 2803 1522 2807
rect 1522 2803 1525 2807
rect 1438 2718 1442 2722
rect 1446 2718 1450 2722
rect 1462 2728 1466 2732
rect 1462 2578 1466 2582
rect 1454 2518 1458 2522
rect 1438 2478 1442 2482
rect 1430 2468 1434 2472
rect 1438 2338 1442 2342
rect 1430 2268 1434 2272
rect 1430 2258 1434 2262
rect 1414 2178 1418 2182
rect 1422 2168 1426 2172
rect 1406 1938 1410 1942
rect 1374 1748 1378 1752
rect 1438 1958 1442 1962
rect 1374 1728 1378 1732
rect 1382 1718 1386 1722
rect 1358 1598 1362 1602
rect 1342 1588 1346 1592
rect 1358 1588 1362 1592
rect 1334 1548 1338 1552
rect 1342 1538 1346 1542
rect 1334 1508 1338 1512
rect 1334 1468 1338 1472
rect 1310 1338 1314 1342
rect 1302 1318 1306 1322
rect 1278 1258 1282 1262
rect 1294 1258 1298 1262
rect 1246 1228 1250 1232
rect 1238 1178 1242 1182
rect 1238 1158 1242 1162
rect 1246 1148 1250 1152
rect 1222 1138 1226 1142
rect 1206 998 1210 1002
rect 1262 1188 1266 1192
rect 1254 1138 1258 1142
rect 1254 1118 1258 1122
rect 1270 1078 1274 1082
rect 1230 1048 1234 1052
rect 1222 988 1226 992
rect 1198 948 1202 952
rect 1206 928 1210 932
rect 1214 918 1218 922
rect 1206 898 1210 902
rect 1198 878 1202 882
rect 1206 858 1210 862
rect 1214 858 1218 862
rect 1206 818 1210 822
rect 1214 818 1218 822
rect 1206 798 1210 802
rect 1254 1018 1258 1022
rect 1246 1008 1250 1012
rect 1254 968 1258 972
rect 1270 1008 1274 1012
rect 1246 938 1250 942
rect 1262 918 1266 922
rect 1262 908 1266 912
rect 1286 1178 1290 1182
rect 1310 1278 1314 1282
rect 1350 1388 1354 1392
rect 1342 1368 1346 1372
rect 1302 1158 1306 1162
rect 1342 1268 1346 1272
rect 1334 1188 1338 1192
rect 1318 1168 1322 1172
rect 1302 1138 1306 1142
rect 1294 1108 1298 1112
rect 1294 1078 1298 1082
rect 1342 1148 1346 1152
rect 1334 1138 1338 1142
rect 1326 1118 1330 1122
rect 1318 1108 1322 1112
rect 1286 1038 1290 1042
rect 1278 968 1282 972
rect 1374 1508 1378 1512
rect 1374 1478 1378 1482
rect 1382 1478 1386 1482
rect 1422 1768 1426 1772
rect 1454 2298 1458 2302
rect 1454 2248 1458 2252
rect 1478 2628 1482 2632
rect 1486 2578 1490 2582
rect 1502 2668 1506 2672
rect 1514 2603 1518 2607
rect 1521 2603 1522 2607
rect 1522 2603 1525 2607
rect 1550 2888 1554 2892
rect 1654 3168 1658 3172
rect 1614 2918 1618 2922
rect 1654 2918 1658 2922
rect 1622 2908 1626 2912
rect 1566 2788 1570 2792
rect 1494 2448 1498 2452
rect 1486 2388 1490 2392
rect 1478 2348 1482 2352
rect 1470 2038 1474 2042
rect 1534 2448 1538 2452
rect 1514 2403 1518 2407
rect 1521 2403 1522 2407
rect 1522 2403 1525 2407
rect 1518 2288 1522 2292
rect 1526 2268 1530 2272
rect 1514 2203 1518 2207
rect 1521 2203 1522 2207
rect 1522 2203 1525 2207
rect 1558 2498 1562 2502
rect 1550 2208 1554 2212
rect 1494 2188 1498 2192
rect 1558 2188 1562 2192
rect 1486 2138 1490 2142
rect 1534 2178 1538 2182
rect 1558 2048 1562 2052
rect 1502 2018 1506 2022
rect 1514 2003 1518 2007
rect 1521 2003 1522 2007
rect 1522 2003 1525 2007
rect 1470 1958 1474 1962
rect 1470 1908 1474 1912
rect 1526 1878 1530 1882
rect 1502 1858 1506 1862
rect 1462 1808 1466 1812
rect 1422 1718 1426 1722
rect 1430 1718 1434 1722
rect 1406 1658 1410 1662
rect 1398 1608 1402 1612
rect 1406 1608 1410 1612
rect 1390 1438 1394 1442
rect 1382 1408 1386 1412
rect 1390 1408 1394 1412
rect 1374 1368 1378 1372
rect 1366 1358 1370 1362
rect 1358 1348 1362 1352
rect 1366 1348 1370 1352
rect 1382 1338 1386 1342
rect 1398 1338 1402 1342
rect 1414 1568 1418 1572
rect 1430 1688 1434 1692
rect 1550 1928 1554 1932
rect 1542 1818 1546 1822
rect 1534 1808 1538 1812
rect 1514 1803 1518 1807
rect 1521 1803 1522 1807
rect 1522 1803 1525 1807
rect 1502 1798 1506 1802
rect 1582 2718 1586 2722
rect 1582 2448 1586 2452
rect 1590 2358 1594 2362
rect 1582 2268 1586 2272
rect 1574 2228 1578 2232
rect 1574 2078 1578 2082
rect 1582 2038 1586 2042
rect 1590 2038 1594 2042
rect 1606 2668 1610 2672
rect 1654 2858 1658 2862
rect 1710 3168 1714 3172
rect 1702 3028 1706 3032
rect 1702 2848 1706 2852
rect 1622 2648 1626 2652
rect 1662 2688 1666 2692
rect 1606 2598 1610 2602
rect 1622 2568 1626 2572
rect 1606 2558 1610 2562
rect 1614 2558 1618 2562
rect 1670 2528 1674 2532
rect 1638 2508 1642 2512
rect 1662 2498 1666 2502
rect 1694 2568 1698 2572
rect 1662 2358 1666 2362
rect 1654 2348 1658 2352
rect 1694 2398 1698 2402
rect 1846 3238 1850 3242
rect 1878 3188 1882 3192
rect 1726 3068 1730 3072
rect 1726 2798 1730 2802
rect 1814 3138 1818 3142
rect 1726 2718 1730 2722
rect 1734 2628 1738 2632
rect 1726 2608 1730 2612
rect 1718 2398 1722 2402
rect 1726 2328 1730 2332
rect 1718 2268 1722 2272
rect 1630 2178 1634 2182
rect 1702 2218 1706 2222
rect 1654 2198 1658 2202
rect 1646 2118 1650 2122
rect 1654 2018 1658 2022
rect 1670 1998 1674 2002
rect 1614 1988 1618 1992
rect 1670 1958 1674 1962
rect 1678 1958 1682 1962
rect 1582 1948 1586 1952
rect 1486 1758 1490 1762
rect 1542 1758 1546 1762
rect 1502 1748 1506 1752
rect 1470 1688 1474 1692
rect 1454 1668 1458 1672
rect 1438 1658 1442 1662
rect 1478 1608 1482 1612
rect 1454 1598 1458 1602
rect 1470 1598 1474 1602
rect 1422 1538 1426 1542
rect 1414 1508 1418 1512
rect 1518 1718 1522 1722
rect 1510 1668 1514 1672
rect 1514 1603 1518 1607
rect 1521 1603 1522 1607
rect 1522 1603 1525 1607
rect 1534 1598 1538 1602
rect 1526 1578 1530 1582
rect 1510 1568 1514 1572
rect 1454 1548 1458 1552
rect 1494 1548 1498 1552
rect 1502 1548 1506 1552
rect 1478 1538 1482 1542
rect 1494 1538 1498 1542
rect 1454 1508 1458 1512
rect 1462 1508 1466 1512
rect 1422 1498 1426 1502
rect 1430 1498 1434 1502
rect 1478 1498 1482 1502
rect 1486 1498 1490 1502
rect 1494 1478 1498 1482
rect 1502 1478 1506 1482
rect 1422 1438 1426 1442
rect 1478 1438 1482 1442
rect 1462 1378 1466 1382
rect 1438 1348 1442 1352
rect 1390 1328 1394 1332
rect 1350 1088 1354 1092
rect 1334 1078 1338 1082
rect 1342 1078 1346 1082
rect 1334 1068 1338 1072
rect 1318 1038 1322 1042
rect 1318 1018 1322 1022
rect 1302 938 1306 942
rect 1310 938 1314 942
rect 1230 878 1234 882
rect 1278 828 1282 832
rect 1294 918 1298 922
rect 1302 908 1306 912
rect 1302 898 1306 902
rect 1294 878 1298 882
rect 1326 988 1330 992
rect 1366 1138 1370 1142
rect 1382 1168 1386 1172
rect 1382 1138 1386 1142
rect 1390 1138 1394 1142
rect 1374 1078 1378 1082
rect 1366 1068 1370 1072
rect 1334 918 1338 922
rect 1342 908 1346 912
rect 1318 898 1322 902
rect 1318 828 1322 832
rect 1286 808 1290 812
rect 1238 788 1242 792
rect 1246 788 1250 792
rect 1246 728 1250 732
rect 1222 718 1226 722
rect 1350 828 1354 832
rect 1326 818 1330 822
rect 1342 768 1346 772
rect 1342 748 1346 752
rect 1350 748 1354 752
rect 1318 738 1322 742
rect 1334 738 1338 742
rect 1422 1258 1426 1262
rect 1430 1258 1434 1262
rect 1422 1238 1426 1242
rect 1406 1158 1410 1162
rect 1430 1188 1434 1192
rect 1574 1788 1578 1792
rect 1646 1928 1650 1932
rect 1622 1918 1626 1922
rect 1630 1918 1634 1922
rect 1598 1898 1602 1902
rect 1598 1858 1602 1862
rect 1630 1858 1634 1862
rect 1590 1818 1594 1822
rect 1582 1738 1586 1742
rect 1566 1698 1570 1702
rect 1614 1798 1618 1802
rect 1606 1788 1610 1792
rect 1598 1718 1602 1722
rect 1558 1668 1562 1672
rect 1550 1608 1554 1612
rect 1590 1668 1594 1672
rect 1566 1578 1570 1582
rect 1518 1458 1522 1462
rect 1542 1458 1546 1462
rect 1558 1478 1562 1482
rect 1582 1568 1586 1572
rect 1574 1558 1578 1562
rect 1638 1788 1642 1792
rect 1670 1918 1674 1922
rect 1654 1848 1658 1852
rect 1654 1788 1658 1792
rect 1686 1878 1690 1882
rect 1702 2038 1706 2042
rect 1782 3048 1786 3052
rect 1814 2938 1818 2942
rect 1790 2928 1794 2932
rect 1766 2918 1770 2922
rect 1758 2698 1762 2702
rect 1750 2398 1754 2402
rect 1742 2348 1746 2352
rect 1750 2328 1754 2332
rect 1782 2848 1786 2852
rect 1798 2768 1802 2772
rect 1790 2738 1794 2742
rect 1774 2568 1778 2572
rect 1766 2558 1770 2562
rect 1782 2558 1786 2562
rect 1742 2158 1746 2162
rect 1726 2058 1730 2062
rect 1734 2058 1738 2062
rect 1734 2038 1738 2042
rect 1726 2028 1730 2032
rect 1758 2098 1762 2102
rect 1782 2378 1786 2382
rect 1782 2358 1786 2362
rect 1774 2348 1778 2352
rect 1790 2208 1794 2212
rect 1774 2168 1778 2172
rect 1766 2038 1770 2042
rect 1718 1928 1722 1932
rect 1694 1868 1698 1872
rect 1734 1868 1738 1872
rect 1742 1868 1746 1872
rect 1710 1858 1714 1862
rect 1718 1858 1722 1862
rect 1862 2988 1866 2992
rect 1862 2918 1866 2922
rect 1878 2908 1882 2912
rect 1846 2888 1850 2892
rect 1846 2858 1850 2862
rect 1870 2768 1874 2772
rect 1838 2618 1842 2622
rect 1894 2878 1898 2882
rect 1926 2928 1930 2932
rect 1926 2808 1930 2812
rect 1862 2578 1866 2582
rect 1838 2528 1842 2532
rect 1846 2528 1850 2532
rect 1854 2518 1858 2522
rect 1830 2328 1834 2332
rect 1830 2288 1834 2292
rect 1846 2198 1850 2202
rect 1846 2148 1850 2152
rect 1798 2128 1802 2132
rect 1790 2118 1794 2122
rect 1782 2018 1786 2022
rect 1774 2008 1778 2012
rect 1782 1928 1786 1932
rect 1798 1928 1802 1932
rect 1766 1898 1770 1902
rect 1790 1908 1794 1912
rect 1774 1888 1778 1892
rect 1758 1878 1762 1882
rect 1702 1848 1706 1852
rect 1750 1848 1754 1852
rect 1686 1808 1690 1812
rect 1662 1688 1666 1692
rect 1654 1678 1658 1682
rect 1630 1588 1634 1592
rect 1614 1578 1618 1582
rect 1590 1548 1594 1552
rect 1598 1548 1602 1552
rect 1534 1438 1538 1442
rect 1510 1428 1514 1432
rect 1502 1418 1506 1422
rect 1494 1408 1498 1412
rect 1534 1408 1538 1412
rect 1514 1403 1518 1407
rect 1521 1403 1522 1407
rect 1522 1403 1525 1407
rect 1478 1288 1482 1292
rect 1486 1288 1490 1292
rect 1470 1268 1474 1272
rect 1446 1238 1450 1242
rect 1438 1168 1442 1172
rect 1422 1118 1426 1122
rect 1454 1188 1458 1192
rect 1462 1148 1466 1152
rect 1494 1208 1498 1212
rect 1514 1203 1518 1207
rect 1521 1203 1522 1207
rect 1522 1203 1525 1207
rect 1502 1198 1506 1202
rect 1486 1128 1490 1132
rect 1470 1118 1474 1122
rect 1478 1088 1482 1092
rect 1486 1088 1490 1092
rect 1454 1078 1458 1082
rect 1438 1058 1442 1062
rect 1414 1008 1418 1012
rect 1366 918 1370 922
rect 1286 728 1290 732
rect 1302 728 1306 732
rect 1254 708 1258 712
rect 1262 708 1266 712
rect 1198 648 1202 652
rect 1214 638 1218 642
rect 1198 628 1202 632
rect 1166 618 1170 622
rect 1174 618 1178 622
rect 1190 618 1194 622
rect 1166 548 1170 552
rect 1182 548 1186 552
rect 1174 538 1178 542
rect 1166 378 1170 382
rect 1158 358 1162 362
rect 1142 348 1146 352
rect 1126 238 1130 242
rect 1142 258 1146 262
rect 1134 168 1138 172
rect 1182 238 1186 242
rect 1174 178 1178 182
rect 1102 118 1106 122
rect 1094 68 1098 72
rect 1142 58 1146 62
rect 1286 668 1290 672
rect 1294 658 1298 662
rect 1270 628 1274 632
rect 1278 598 1282 602
rect 1294 558 1298 562
rect 1278 538 1282 542
rect 1334 668 1338 672
rect 1310 608 1314 612
rect 1318 608 1322 612
rect 1318 568 1322 572
rect 1334 568 1338 572
rect 1310 558 1314 562
rect 1302 548 1306 552
rect 1310 548 1314 552
rect 1326 538 1330 542
rect 1294 528 1298 532
rect 1254 428 1258 432
rect 1262 428 1266 432
rect 1230 408 1234 412
rect 1182 78 1186 82
rect 1214 358 1218 362
rect 1270 378 1274 382
rect 1222 218 1226 222
rect 1110 28 1114 32
rect 1230 58 1234 62
rect 1270 228 1274 232
rect 1254 188 1258 192
rect 1246 88 1250 92
rect 1230 48 1234 52
rect 1286 88 1290 92
rect 1334 518 1338 522
rect 1422 988 1426 992
rect 1438 988 1442 992
rect 1406 958 1410 962
rect 1390 888 1394 892
rect 1406 928 1410 932
rect 1422 888 1426 892
rect 1374 848 1378 852
rect 1398 848 1402 852
rect 1438 848 1442 852
rect 1406 808 1410 812
rect 1390 698 1394 702
rect 1462 1068 1466 1072
rect 1462 1038 1466 1042
rect 1470 1038 1474 1042
rect 1542 1298 1546 1302
rect 1566 1398 1570 1402
rect 1558 1368 1562 1372
rect 1630 1548 1634 1552
rect 1654 1558 1658 1562
rect 1606 1488 1610 1492
rect 1590 1478 1594 1482
rect 1630 1478 1634 1482
rect 1614 1468 1618 1472
rect 1606 1438 1610 1442
rect 1614 1428 1618 1432
rect 1550 1288 1554 1292
rect 1566 1288 1570 1292
rect 1542 1268 1546 1272
rect 1582 1338 1586 1342
rect 1598 1358 1602 1362
rect 1654 1478 1658 1482
rect 1654 1438 1658 1442
rect 1606 1338 1610 1342
rect 1550 1248 1554 1252
rect 1550 1208 1554 1212
rect 1542 1168 1546 1172
rect 1542 1138 1546 1142
rect 1526 1048 1530 1052
rect 1534 1048 1538 1052
rect 1502 1008 1506 1012
rect 1486 978 1490 982
rect 1430 738 1434 742
rect 1406 728 1410 732
rect 1390 578 1394 582
rect 1390 518 1394 522
rect 1326 288 1330 292
rect 1310 268 1314 272
rect 1310 238 1314 242
rect 1302 98 1306 102
rect 1334 158 1338 162
rect 1318 138 1322 142
rect 1342 108 1346 112
rect 1406 638 1410 642
rect 1406 538 1410 542
rect 1406 518 1410 522
rect 1470 898 1474 902
rect 1514 1003 1518 1007
rect 1521 1003 1522 1007
rect 1522 1003 1525 1007
rect 1502 998 1506 1002
rect 1502 928 1506 932
rect 1494 918 1498 922
rect 1502 868 1506 872
rect 1478 858 1482 862
rect 1478 778 1482 782
rect 1510 828 1514 832
rect 1514 803 1518 807
rect 1521 803 1522 807
rect 1522 803 1525 807
rect 1502 798 1506 802
rect 1462 758 1466 762
rect 1486 758 1490 762
rect 1566 1198 1570 1202
rect 1590 1208 1594 1212
rect 1558 1078 1562 1082
rect 1550 968 1554 972
rect 1558 918 1562 922
rect 1574 1138 1578 1142
rect 1598 1148 1602 1152
rect 1622 1228 1626 1232
rect 1638 1268 1642 1272
rect 1622 1138 1626 1142
rect 1614 1128 1618 1132
rect 1598 1108 1602 1112
rect 1622 1088 1626 1092
rect 1614 1068 1618 1072
rect 1582 1008 1586 1012
rect 1590 1008 1594 1012
rect 1590 958 1594 962
rect 1598 958 1602 962
rect 1558 798 1562 802
rect 1518 788 1522 792
rect 1542 738 1546 742
rect 1494 728 1498 732
rect 1470 708 1474 712
rect 1454 668 1458 672
rect 1438 658 1442 662
rect 1422 628 1426 632
rect 1422 548 1426 552
rect 1414 488 1418 492
rect 1422 488 1426 492
rect 1422 458 1426 462
rect 1486 658 1490 662
rect 1470 628 1474 632
rect 1486 618 1490 622
rect 1486 598 1490 602
rect 1518 698 1522 702
rect 1526 688 1530 692
rect 1510 678 1514 682
rect 1502 668 1506 672
rect 1614 908 1618 912
rect 1678 1698 1682 1702
rect 1758 1838 1762 1842
rect 1710 1818 1714 1822
rect 1750 1818 1754 1822
rect 1718 1788 1722 1792
rect 1702 1768 1706 1772
rect 1694 1698 1698 1702
rect 1774 1808 1778 1812
rect 1790 1748 1794 1752
rect 1798 1718 1802 1722
rect 1718 1648 1722 1652
rect 1726 1648 1730 1652
rect 1710 1608 1714 1612
rect 1694 1598 1698 1602
rect 1686 1588 1690 1592
rect 1678 1578 1682 1582
rect 1686 1568 1690 1572
rect 1710 1588 1714 1592
rect 1710 1568 1714 1572
rect 1678 1498 1682 1502
rect 1766 1698 1770 1702
rect 1790 1688 1794 1692
rect 1798 1688 1802 1692
rect 1766 1668 1770 1672
rect 1766 1618 1770 1622
rect 1750 1578 1754 1582
rect 1734 1558 1738 1562
rect 1734 1438 1738 1442
rect 1790 1608 1794 1612
rect 1766 1598 1770 1602
rect 1774 1558 1778 1562
rect 1766 1548 1770 1552
rect 1766 1478 1770 1482
rect 1774 1478 1778 1482
rect 1774 1438 1778 1442
rect 1766 1428 1770 1432
rect 1782 1428 1786 1432
rect 1750 1408 1754 1412
rect 1758 1408 1762 1412
rect 1702 1398 1706 1402
rect 1750 1398 1754 1402
rect 1758 1398 1762 1402
rect 1694 1358 1698 1362
rect 1678 1338 1682 1342
rect 1670 1228 1674 1232
rect 1646 1198 1650 1202
rect 1630 1038 1634 1042
rect 1646 1038 1650 1042
rect 1630 968 1634 972
rect 1638 848 1642 852
rect 1598 748 1602 752
rect 1582 698 1586 702
rect 1574 688 1578 692
rect 1502 608 1506 612
rect 1550 608 1554 612
rect 1514 603 1518 607
rect 1521 603 1522 607
rect 1522 603 1525 607
rect 1494 478 1498 482
rect 1454 468 1458 472
rect 1438 398 1442 402
rect 1514 403 1518 407
rect 1521 403 1522 407
rect 1522 403 1525 407
rect 1422 308 1426 312
rect 1478 288 1482 292
rect 1430 278 1434 282
rect 1470 278 1474 282
rect 1390 148 1394 152
rect 1438 148 1442 152
rect 1374 98 1378 102
rect 1350 88 1354 92
rect 1350 58 1354 62
rect 1430 88 1434 92
rect 1438 58 1442 62
rect 1478 108 1482 112
rect 1470 48 1474 52
rect 1566 458 1570 462
rect 1614 698 1618 702
rect 1662 1118 1666 1122
rect 1670 1108 1674 1112
rect 1670 1068 1674 1072
rect 1670 1018 1674 1022
rect 1662 998 1666 1002
rect 1622 568 1626 572
rect 1590 428 1594 432
rect 1614 428 1618 432
rect 1598 278 1602 282
rect 1574 258 1578 262
rect 1514 203 1518 207
rect 1521 203 1522 207
rect 1522 203 1525 207
rect 1502 128 1506 132
rect 1494 78 1498 82
rect 1694 1338 1698 1342
rect 1686 1328 1690 1332
rect 1766 1338 1770 1342
rect 1750 1328 1754 1332
rect 1766 1328 1770 1332
rect 1718 1318 1722 1322
rect 1702 1298 1706 1302
rect 1718 1298 1722 1302
rect 1702 1228 1706 1232
rect 1710 1228 1714 1232
rect 1694 1208 1698 1212
rect 1686 1128 1690 1132
rect 1702 1158 1706 1162
rect 1734 1308 1738 1312
rect 1750 1308 1754 1312
rect 1758 1288 1762 1292
rect 1726 1198 1730 1202
rect 1790 1398 1794 1402
rect 1782 1298 1786 1302
rect 1782 1278 1786 1282
rect 1846 2118 1850 2122
rect 1878 2378 1882 2382
rect 1870 2368 1874 2372
rect 1894 2568 1898 2572
rect 1902 2558 1906 2562
rect 1918 2608 1922 2612
rect 1862 2318 1866 2322
rect 1910 2318 1914 2322
rect 1894 2308 1898 2312
rect 1894 2178 1898 2182
rect 1926 2138 1930 2142
rect 1918 2088 1922 2092
rect 1902 2058 1906 2062
rect 1862 2048 1866 2052
rect 1830 2028 1834 2032
rect 1830 2008 1834 2012
rect 1838 1998 1842 2002
rect 1846 1988 1850 1992
rect 1854 1958 1858 1962
rect 1854 1938 1858 1942
rect 1830 1918 1834 1922
rect 1830 1898 1834 1902
rect 1910 2048 1914 2052
rect 1926 2028 1930 2032
rect 1942 2858 1946 2862
rect 1990 3128 1994 3132
rect 1982 3048 1986 3052
rect 1966 2738 1970 2742
rect 1990 2868 1994 2872
rect 2166 3288 2170 3292
rect 2182 3268 2186 3272
rect 2030 3258 2034 3262
rect 2026 3103 2030 3107
rect 2033 3103 2034 3107
rect 2034 3103 2037 3107
rect 2006 3088 2010 3092
rect 2166 3128 2170 3132
rect 2054 2948 2058 2952
rect 2022 2938 2026 2942
rect 1990 2858 1994 2862
rect 1998 2728 2002 2732
rect 2006 2708 2010 2712
rect 2026 2903 2030 2907
rect 2033 2903 2034 2907
rect 2034 2903 2037 2907
rect 2102 3068 2106 3072
rect 2086 2918 2090 2922
rect 2078 2888 2082 2892
rect 2070 2748 2074 2752
rect 2062 2728 2066 2732
rect 2026 2703 2030 2707
rect 2033 2703 2034 2707
rect 2034 2703 2037 2707
rect 2014 2698 2018 2702
rect 2006 2608 2010 2612
rect 1950 2358 1954 2362
rect 1966 2358 1970 2362
rect 1942 2328 1946 2332
rect 1950 2318 1954 2322
rect 1958 2318 1962 2322
rect 1878 1958 1882 1962
rect 1854 1848 1858 1852
rect 1838 1798 1842 1802
rect 1814 1718 1818 1722
rect 1846 1768 1850 1772
rect 1862 1838 1866 1842
rect 1870 1838 1874 1842
rect 1886 1908 1890 1912
rect 1918 1918 1922 1922
rect 1894 1888 1898 1892
rect 1902 1868 1906 1872
rect 1862 1768 1866 1772
rect 1846 1728 1850 1732
rect 1822 1668 1826 1672
rect 1806 1548 1810 1552
rect 1814 1448 1818 1452
rect 1830 1448 1834 1452
rect 1822 1368 1826 1372
rect 1806 1338 1810 1342
rect 1798 1298 1802 1302
rect 1782 1228 1786 1232
rect 1758 1198 1762 1202
rect 1742 1188 1746 1192
rect 1750 1188 1754 1192
rect 1734 1158 1738 1162
rect 1742 1158 1746 1162
rect 1718 1118 1722 1122
rect 1702 1098 1706 1102
rect 1694 1088 1698 1092
rect 1718 1078 1722 1082
rect 1686 1018 1690 1022
rect 1694 1008 1698 1012
rect 1678 958 1682 962
rect 1670 908 1674 912
rect 1670 778 1674 782
rect 1734 1068 1738 1072
rect 1750 1038 1754 1042
rect 1726 948 1730 952
rect 1734 948 1738 952
rect 1774 1168 1778 1172
rect 1702 918 1706 922
rect 1718 918 1722 922
rect 1702 878 1706 882
rect 1686 798 1690 802
rect 1694 798 1698 802
rect 1742 908 1746 912
rect 1750 898 1754 902
rect 1726 878 1730 882
rect 1758 798 1762 802
rect 1686 778 1690 782
rect 1766 778 1770 782
rect 1822 1348 1826 1352
rect 1822 1298 1826 1302
rect 1846 1408 1850 1412
rect 1846 1368 1850 1372
rect 1846 1358 1850 1362
rect 1894 1838 1898 1842
rect 1878 1678 1882 1682
rect 1886 1678 1890 1682
rect 1862 1588 1866 1592
rect 1870 1578 1874 1582
rect 1862 1548 1866 1552
rect 1910 1838 1914 1842
rect 2014 2598 2018 2602
rect 2038 2528 2042 2532
rect 2026 2503 2030 2507
rect 2033 2503 2034 2507
rect 2034 2503 2037 2507
rect 2006 2308 2010 2312
rect 2026 2303 2030 2307
rect 2033 2303 2034 2307
rect 2034 2303 2037 2307
rect 2046 2298 2050 2302
rect 2022 2278 2026 2282
rect 2062 2518 2066 2522
rect 2070 2498 2074 2502
rect 2070 2338 2074 2342
rect 2070 2258 2074 2262
rect 2110 2868 2114 2872
rect 2126 2718 2130 2722
rect 2102 2668 2106 2672
rect 2142 2638 2146 2642
rect 2134 2568 2138 2572
rect 2182 3068 2186 3072
rect 2238 3288 2242 3292
rect 2214 3248 2218 3252
rect 2222 3138 2226 3142
rect 2206 3098 2210 3102
rect 2182 2948 2186 2952
rect 2206 2858 2210 2862
rect 2134 2488 2138 2492
rect 2118 2358 2122 2362
rect 2102 2348 2106 2352
rect 2102 2318 2106 2322
rect 2102 2288 2106 2292
rect 2094 2268 2098 2272
rect 2086 2218 2090 2222
rect 2062 2178 2066 2182
rect 2142 2278 2146 2282
rect 2110 2268 2114 2272
rect 2126 2248 2130 2252
rect 1958 2148 1962 2152
rect 2046 2128 2050 2132
rect 2026 2103 2030 2107
rect 2033 2103 2034 2107
rect 2034 2103 2037 2107
rect 2054 2098 2058 2102
rect 2134 2118 2138 2122
rect 2134 2098 2138 2102
rect 2062 2058 2066 2062
rect 1942 1948 1946 1952
rect 1950 1898 1954 1902
rect 1942 1868 1946 1872
rect 1934 1798 1938 1802
rect 1934 1778 1938 1782
rect 1926 1768 1930 1772
rect 1910 1758 1914 1762
rect 1942 1768 1946 1772
rect 1926 1728 1930 1732
rect 1918 1678 1922 1682
rect 1902 1598 1906 1602
rect 1886 1558 1890 1562
rect 1886 1538 1890 1542
rect 1894 1538 1898 1542
rect 1894 1498 1898 1502
rect 1878 1488 1882 1492
rect 1886 1488 1890 1492
rect 1894 1398 1898 1402
rect 1870 1388 1874 1392
rect 1894 1378 1898 1382
rect 1870 1358 1874 1362
rect 1894 1358 1898 1362
rect 1878 1348 1882 1352
rect 1878 1328 1882 1332
rect 1886 1328 1890 1332
rect 1862 1318 1866 1322
rect 1878 1318 1882 1322
rect 1838 1218 1842 1222
rect 1830 1208 1834 1212
rect 1838 1208 1842 1212
rect 1814 1178 1818 1182
rect 1798 1138 1802 1142
rect 1814 1138 1818 1142
rect 1790 1128 1794 1132
rect 1806 1128 1810 1132
rect 1806 1108 1810 1112
rect 1806 1088 1810 1092
rect 1814 1088 1818 1092
rect 1782 848 1786 852
rect 1718 748 1722 752
rect 1734 748 1738 752
rect 1798 898 1802 902
rect 1798 888 1802 892
rect 1830 1108 1834 1112
rect 1870 1218 1874 1222
rect 1902 1318 1906 1322
rect 1974 1968 1978 1972
rect 1990 1968 1994 1972
rect 2038 1928 2042 1932
rect 1998 1918 2002 1922
rect 2126 2048 2130 2052
rect 2198 2568 2202 2572
rect 2190 2548 2194 2552
rect 2174 2528 2178 2532
rect 2310 3268 2314 3272
rect 2374 3108 2378 3112
rect 2310 3048 2314 3052
rect 2438 3068 2442 3072
rect 2382 3058 2386 3062
rect 2246 2868 2250 2872
rect 2246 2668 2250 2672
rect 2214 2628 2218 2632
rect 2206 2558 2210 2562
rect 2206 2518 2210 2522
rect 2166 2288 2170 2292
rect 2166 2278 2170 2282
rect 2198 2268 2202 2272
rect 2206 2258 2210 2262
rect 2174 2248 2178 2252
rect 2182 2168 2186 2172
rect 2222 2618 2226 2622
rect 2166 2088 2170 2092
rect 2206 2088 2210 2092
rect 2230 2368 2234 2372
rect 2150 2048 2154 2052
rect 2110 1998 2114 2002
rect 2062 1958 2066 1962
rect 2086 1958 2090 1962
rect 2014 1908 2018 1912
rect 2026 1903 2030 1907
rect 2033 1903 2034 1907
rect 2034 1903 2037 1907
rect 1990 1858 1994 1862
rect 2014 1858 2018 1862
rect 2022 1858 2026 1862
rect 1998 1838 2002 1842
rect 2038 1838 2042 1842
rect 2022 1828 2026 1832
rect 1998 1798 2002 1802
rect 1982 1728 1986 1732
rect 1958 1698 1962 1702
rect 2038 1768 2042 1772
rect 2014 1708 2018 1712
rect 1942 1688 1946 1692
rect 1934 1548 1938 1552
rect 1958 1668 1962 1672
rect 1982 1658 1986 1662
rect 1950 1588 1954 1592
rect 1966 1588 1970 1592
rect 1958 1578 1962 1582
rect 1926 1498 1930 1502
rect 1934 1498 1938 1502
rect 1942 1428 1946 1432
rect 1942 1358 1946 1362
rect 1926 1348 1930 1352
rect 1934 1348 1938 1352
rect 1918 1298 1922 1302
rect 1902 1288 1906 1292
rect 1902 1258 1906 1262
rect 1894 1188 1898 1192
rect 1846 1098 1850 1102
rect 1822 1058 1826 1062
rect 1838 958 1842 962
rect 1846 958 1850 962
rect 1862 978 1866 982
rect 1878 1128 1882 1132
rect 1886 1128 1890 1132
rect 1878 1108 1882 1112
rect 1830 928 1834 932
rect 1862 858 1866 862
rect 1830 848 1834 852
rect 1846 848 1850 852
rect 1894 1078 1898 1082
rect 1910 1058 1914 1062
rect 1902 1038 1906 1042
rect 1886 938 1890 942
rect 1878 918 1882 922
rect 1870 818 1874 822
rect 1790 798 1794 802
rect 1846 748 1850 752
rect 1854 738 1858 742
rect 1790 708 1794 712
rect 1782 698 1786 702
rect 1710 658 1714 662
rect 1782 678 1786 682
rect 1766 668 1770 672
rect 1790 658 1794 662
rect 1702 648 1706 652
rect 1734 648 1738 652
rect 1718 528 1722 532
rect 1742 478 1746 482
rect 1774 458 1778 462
rect 1654 438 1658 442
rect 1678 278 1682 282
rect 1702 348 1706 352
rect 1774 348 1778 352
rect 1686 268 1690 272
rect 1702 268 1706 272
rect 1758 268 1762 272
rect 1766 258 1770 262
rect 1822 688 1826 692
rect 1814 678 1818 682
rect 1822 658 1826 662
rect 1814 558 1818 562
rect 1798 508 1802 512
rect 1854 648 1858 652
rect 1870 698 1874 702
rect 1942 1308 1946 1312
rect 1942 1288 1946 1292
rect 1950 1258 1954 1262
rect 1950 1178 1954 1182
rect 1934 1148 1938 1152
rect 1934 1108 1938 1112
rect 1926 1058 1930 1062
rect 2026 1703 2030 1707
rect 2033 1703 2034 1707
rect 2034 1703 2037 1707
rect 2102 1948 2106 1952
rect 2070 1828 2074 1832
rect 2062 1728 2066 1732
rect 2054 1708 2058 1712
rect 2046 1648 2050 1652
rect 2086 1808 2090 1812
rect 2086 1788 2090 1792
rect 2110 1928 2114 1932
rect 2126 1918 2130 1922
rect 2110 1858 2114 1862
rect 2118 1858 2122 1862
rect 2094 1778 2098 1782
rect 2118 1768 2122 1772
rect 2086 1748 2090 1752
rect 2182 2058 2186 2062
rect 2262 2528 2266 2532
rect 2366 2928 2370 2932
rect 2310 2668 2314 2672
rect 2254 2178 2258 2182
rect 2278 2498 2282 2502
rect 2270 2328 2274 2332
rect 2270 2288 2274 2292
rect 2198 1978 2202 1982
rect 2158 1908 2162 1912
rect 2142 1818 2146 1822
rect 2134 1748 2138 1752
rect 2118 1718 2122 1722
rect 2078 1678 2082 1682
rect 2110 1678 2114 1682
rect 2062 1598 2066 1602
rect 2054 1588 2058 1592
rect 2014 1578 2018 1582
rect 1966 1568 1970 1572
rect 2006 1568 2010 1572
rect 1990 1558 1994 1562
rect 2006 1558 2010 1562
rect 2046 1558 2050 1562
rect 1974 1548 1978 1552
rect 1966 1378 1970 1382
rect 1982 1538 1986 1542
rect 2094 1588 2098 1592
rect 2070 1548 2074 1552
rect 2006 1508 2010 1512
rect 2026 1503 2030 1507
rect 2033 1503 2034 1507
rect 2034 1503 2037 1507
rect 2118 1618 2122 1622
rect 2110 1578 2114 1582
rect 2118 1558 2122 1562
rect 2054 1538 2058 1542
rect 2006 1498 2010 1502
rect 2046 1498 2050 1502
rect 1990 1488 1994 1492
rect 2038 1468 2042 1472
rect 1998 1428 2002 1432
rect 1990 1368 1994 1372
rect 1982 1318 1986 1322
rect 1974 1298 1978 1302
rect 1974 1218 1978 1222
rect 1982 1218 1986 1222
rect 1966 1168 1970 1172
rect 1958 1128 1962 1132
rect 1958 1108 1962 1112
rect 1966 1108 1970 1112
rect 2030 1418 2034 1422
rect 2014 1358 2018 1362
rect 2006 1328 2010 1332
rect 2030 1348 2034 1352
rect 2102 1528 2106 1532
rect 2118 1528 2122 1532
rect 2054 1428 2058 1432
rect 2054 1408 2058 1412
rect 2062 1408 2066 1412
rect 2046 1328 2050 1332
rect 2046 1308 2050 1312
rect 2054 1308 2058 1312
rect 2026 1303 2030 1307
rect 2033 1303 2034 1307
rect 2034 1303 2037 1307
rect 2006 1168 2010 1172
rect 1982 1148 1986 1152
rect 1990 1118 1994 1122
rect 1934 1038 1938 1042
rect 1958 1038 1962 1042
rect 1902 978 1906 982
rect 1926 948 1930 952
rect 1958 948 1962 952
rect 1974 948 1978 952
rect 1942 938 1946 942
rect 1950 938 1954 942
rect 1966 918 1970 922
rect 1950 898 1954 902
rect 2006 1098 2010 1102
rect 1998 978 2002 982
rect 1942 878 1946 882
rect 1926 868 1930 872
rect 1966 868 1970 872
rect 1934 848 1938 852
rect 1918 828 1922 832
rect 1910 818 1914 822
rect 1846 618 1850 622
rect 1878 618 1882 622
rect 1830 498 1834 502
rect 1838 348 1842 352
rect 1806 288 1810 292
rect 1838 308 1842 312
rect 1830 288 1834 292
rect 1902 778 1906 782
rect 1934 748 1938 752
rect 1894 598 1898 602
rect 1862 388 1866 392
rect 1934 648 1938 652
rect 1918 618 1922 622
rect 1990 828 1994 832
rect 1990 758 1994 762
rect 1950 738 1954 742
rect 1966 738 1970 742
rect 1950 608 1954 612
rect 1918 438 1922 442
rect 1918 428 1922 432
rect 1814 278 1818 282
rect 1862 278 1866 282
rect 1806 268 1810 272
rect 1822 238 1826 242
rect 1966 538 1970 542
rect 2054 1258 2058 1262
rect 2038 1218 2042 1222
rect 2078 1418 2082 1422
rect 2102 1498 2106 1502
rect 2086 1378 2090 1382
rect 2118 1468 2122 1472
rect 2110 1418 2114 1422
rect 2102 1368 2106 1372
rect 2078 1348 2082 1352
rect 2086 1348 2090 1352
rect 2070 1198 2074 1202
rect 2094 1328 2098 1332
rect 2110 1328 2114 1332
rect 2094 1318 2098 1322
rect 2102 1298 2106 1302
rect 2094 1258 2098 1262
rect 2062 1148 2066 1152
rect 2070 1148 2074 1152
rect 2026 1103 2030 1107
rect 2033 1103 2034 1107
rect 2034 1103 2037 1107
rect 2022 1028 2026 1032
rect 2046 998 2050 1002
rect 2022 958 2026 962
rect 2014 918 2018 922
rect 2026 903 2030 907
rect 2033 903 2034 907
rect 2034 903 2037 907
rect 2014 888 2018 892
rect 2022 888 2026 892
rect 2078 1128 2082 1132
rect 2062 1108 2066 1112
rect 2070 1048 2074 1052
rect 2062 1028 2066 1032
rect 2062 948 2066 952
rect 2038 848 2042 852
rect 2030 818 2034 822
rect 2046 818 2050 822
rect 2070 908 2074 912
rect 2070 868 2074 872
rect 2062 788 2066 792
rect 2062 768 2066 772
rect 2014 738 2018 742
rect 2054 738 2058 742
rect 2014 728 2018 732
rect 2070 708 2074 712
rect 2026 703 2030 707
rect 2033 703 2034 707
rect 2034 703 2037 707
rect 2070 658 2074 662
rect 2086 1108 2090 1112
rect 2094 1048 2098 1052
rect 2086 898 2090 902
rect 2086 858 2090 862
rect 2190 1838 2194 1842
rect 2198 1778 2202 1782
rect 2166 1758 2170 1762
rect 2190 1648 2194 1652
rect 2182 1598 2186 1602
rect 2150 1578 2154 1582
rect 2150 1568 2154 1572
rect 2134 1558 2138 1562
rect 2166 1558 2170 1562
rect 2158 1518 2162 1522
rect 2134 1418 2138 1422
rect 2118 1308 2122 1312
rect 2118 1248 2122 1252
rect 2174 1508 2178 1512
rect 2230 1908 2234 1912
rect 2214 1898 2218 1902
rect 2286 2458 2290 2462
rect 2310 2388 2314 2392
rect 2286 2068 2290 2072
rect 2294 2038 2298 2042
rect 2222 1888 2226 1892
rect 2238 1888 2242 1892
rect 2278 1868 2282 1872
rect 2278 1848 2282 1852
rect 2230 1798 2234 1802
rect 2214 1778 2218 1782
rect 2222 1728 2226 1732
rect 2214 1688 2218 1692
rect 2214 1618 2218 1622
rect 2206 1558 2210 1562
rect 2222 1538 2226 1542
rect 2206 1498 2210 1502
rect 2198 1448 2202 1452
rect 2262 1768 2266 1772
rect 2238 1728 2242 1732
rect 2246 1598 2250 1602
rect 2230 1508 2234 1512
rect 2214 1438 2218 1442
rect 2246 1538 2250 1542
rect 2246 1498 2250 1502
rect 2270 1648 2274 1652
rect 2350 2498 2354 2502
rect 2350 2448 2354 2452
rect 2350 2398 2354 2402
rect 2334 2358 2338 2362
rect 2342 2058 2346 2062
rect 2302 1948 2306 1952
rect 2302 1858 2306 1862
rect 2326 1908 2330 1912
rect 2334 1838 2338 1842
rect 2334 1708 2338 1712
rect 2302 1558 2306 1562
rect 2278 1548 2282 1552
rect 2286 1548 2290 1552
rect 2270 1518 2274 1522
rect 2262 1468 2266 1472
rect 2302 1538 2306 1542
rect 2286 1518 2290 1522
rect 2318 1618 2322 1622
rect 2318 1598 2322 1602
rect 2334 1608 2338 1612
rect 2326 1578 2330 1582
rect 2334 1578 2338 1582
rect 2374 2768 2378 2772
rect 2366 2658 2370 2662
rect 2366 2648 2370 2652
rect 2390 2888 2394 2892
rect 2382 2268 2386 2272
rect 2382 2078 2386 2082
rect 2398 2668 2402 2672
rect 2414 2648 2418 2652
rect 2406 2628 2410 2632
rect 2406 2588 2410 2592
rect 2430 2578 2434 2582
rect 2438 2508 2442 2512
rect 2438 2408 2442 2412
rect 2510 3248 2514 3252
rect 2494 3158 2498 3162
rect 2502 3068 2506 3072
rect 2502 3058 2506 3062
rect 2478 2858 2482 2862
rect 2494 2668 2498 2672
rect 2502 2648 2506 2652
rect 2510 2588 2514 2592
rect 2486 2518 2490 2522
rect 2470 2458 2474 2462
rect 2538 3203 2542 3207
rect 2545 3203 2546 3207
rect 2546 3203 2549 3207
rect 2558 3018 2562 3022
rect 2538 3003 2542 3007
rect 2545 3003 2546 3007
rect 2546 3003 2549 3007
rect 2558 2858 2562 2862
rect 2582 2818 2586 2822
rect 2538 2803 2542 2807
rect 2545 2803 2546 2807
rect 2546 2803 2549 2807
rect 2558 2758 2562 2762
rect 2538 2603 2542 2607
rect 2545 2603 2546 2607
rect 2546 2603 2549 2607
rect 2526 2528 2530 2532
rect 2542 2458 2546 2462
rect 2382 1918 2386 1922
rect 2358 1728 2362 1732
rect 2350 1688 2354 1692
rect 2318 1528 2322 1532
rect 2302 1478 2306 1482
rect 2302 1458 2306 1462
rect 2270 1448 2274 1452
rect 2230 1398 2234 1402
rect 2222 1378 2226 1382
rect 2182 1348 2186 1352
rect 2182 1328 2186 1332
rect 2166 1298 2170 1302
rect 2158 1288 2162 1292
rect 2150 1268 2154 1272
rect 2142 1248 2146 1252
rect 2142 1158 2146 1162
rect 2126 1078 2130 1082
rect 2182 1278 2186 1282
rect 2174 1178 2178 1182
rect 2230 1368 2234 1372
rect 2238 1368 2242 1372
rect 2222 1358 2226 1362
rect 2206 1228 2210 1232
rect 2190 1208 2194 1212
rect 2182 1168 2186 1172
rect 2174 1138 2178 1142
rect 2166 1088 2170 1092
rect 2174 1088 2178 1092
rect 2134 1058 2138 1062
rect 2158 1058 2162 1062
rect 2174 1038 2178 1042
rect 2190 1038 2194 1042
rect 2118 958 2122 962
rect 2174 958 2178 962
rect 2102 898 2106 902
rect 2158 898 2162 902
rect 2118 768 2122 772
rect 2086 678 2090 682
rect 2150 808 2154 812
rect 2142 798 2146 802
rect 2142 758 2146 762
rect 2158 738 2162 742
rect 1998 648 2002 652
rect 2078 648 2082 652
rect 1934 508 1938 512
rect 1958 368 1962 372
rect 1942 308 1946 312
rect 2086 598 2090 602
rect 2026 503 2030 507
rect 2033 503 2034 507
rect 2034 503 2037 507
rect 2150 668 2154 672
rect 2174 888 2178 892
rect 2182 808 2186 812
rect 2182 788 2186 792
rect 2166 608 2170 612
rect 2174 478 2178 482
rect 2006 438 2010 442
rect 2006 328 2010 332
rect 2118 328 2122 332
rect 2014 318 2018 322
rect 2026 303 2030 307
rect 2033 303 2034 307
rect 2034 303 2037 307
rect 1974 268 1978 272
rect 1982 238 1986 242
rect 1798 148 1802 152
rect 1982 178 1986 182
rect 1806 138 1810 142
rect 1798 128 1802 132
rect 1710 108 1714 112
rect 1798 78 1802 82
rect 1622 58 1626 62
rect 1886 98 1890 102
rect 1918 78 1922 82
rect 1974 78 1978 82
rect 2062 268 2066 272
rect 2086 258 2090 262
rect 2062 158 2066 162
rect 2094 158 2098 162
rect 2118 158 2122 162
rect 2026 103 2030 107
rect 2033 103 2034 107
rect 2034 103 2037 107
rect 2158 308 2162 312
rect 2246 1308 2250 1312
rect 2230 1238 2234 1242
rect 2230 1128 2234 1132
rect 2206 1068 2210 1072
rect 2222 1028 2226 1032
rect 2270 1358 2274 1362
rect 2278 1358 2282 1362
rect 2262 1348 2266 1352
rect 2262 1258 2266 1262
rect 2270 1168 2274 1172
rect 2254 1088 2258 1092
rect 2246 1078 2250 1082
rect 2230 958 2234 962
rect 2214 928 2218 932
rect 2206 878 2210 882
rect 2238 868 2242 872
rect 2206 808 2210 812
rect 2198 728 2202 732
rect 2230 768 2234 772
rect 2286 1278 2290 1282
rect 2286 1258 2290 1262
rect 2302 1328 2306 1332
rect 2302 1238 2306 1242
rect 2294 1138 2298 1142
rect 2310 1118 2314 1122
rect 2294 1088 2298 1092
rect 2262 998 2266 1002
rect 2270 998 2274 1002
rect 2278 978 2282 982
rect 2286 978 2290 982
rect 2262 868 2266 872
rect 2302 938 2306 942
rect 2310 868 2314 872
rect 2278 748 2282 752
rect 2278 738 2282 742
rect 2294 718 2298 722
rect 2254 628 2258 632
rect 2134 268 2138 272
rect 2166 238 2170 242
rect 2142 148 2146 152
rect 2182 148 2186 152
rect 2142 108 2146 112
rect 2014 98 2018 102
rect 2062 78 2066 82
rect 2006 68 2010 72
rect 2214 318 2218 322
rect 2238 258 2242 262
rect 2222 68 2226 72
rect 2334 1498 2338 1502
rect 2342 1488 2346 1492
rect 2374 1678 2378 1682
rect 2358 1618 2362 1622
rect 2366 1618 2370 1622
rect 2358 1598 2362 1602
rect 2358 1568 2362 1572
rect 2358 1498 2362 1502
rect 2358 1428 2362 1432
rect 2358 1398 2362 1402
rect 2350 1358 2354 1362
rect 2366 1368 2370 1372
rect 2350 1278 2354 1282
rect 2358 1278 2362 1282
rect 2334 1228 2338 1232
rect 2350 1218 2354 1222
rect 2358 1218 2362 1222
rect 2326 1028 2330 1032
rect 2350 1128 2354 1132
rect 2350 1118 2354 1122
rect 2350 1078 2354 1082
rect 2350 948 2354 952
rect 2334 768 2338 772
rect 2302 618 2306 622
rect 2502 2328 2506 2332
rect 2422 2078 2426 2082
rect 2422 2048 2426 2052
rect 2438 1928 2442 1932
rect 2430 1878 2434 1882
rect 2406 1858 2410 1862
rect 2422 1758 2426 1762
rect 2406 1728 2410 1732
rect 2398 1718 2402 1722
rect 2430 1718 2434 1722
rect 2438 1628 2442 1632
rect 2406 1618 2410 1622
rect 2422 1578 2426 1582
rect 2526 2418 2530 2422
rect 2538 2403 2542 2407
rect 2545 2403 2546 2407
rect 2546 2403 2549 2407
rect 2590 2658 2594 2662
rect 2590 2558 2594 2562
rect 2766 3258 2770 3262
rect 2702 3158 2706 3162
rect 2782 3148 2786 3152
rect 2766 3138 2770 3142
rect 2614 2578 2618 2582
rect 2598 2338 2602 2342
rect 2598 2318 2602 2322
rect 2574 2278 2578 2282
rect 2566 2228 2570 2232
rect 2518 2208 2522 2212
rect 2538 2203 2542 2207
rect 2545 2203 2546 2207
rect 2546 2203 2549 2207
rect 2526 2138 2530 2142
rect 2526 2118 2530 2122
rect 2598 2268 2602 2272
rect 2582 2108 2586 2112
rect 2486 2048 2490 2052
rect 2526 2008 2530 2012
rect 2502 1938 2506 1942
rect 2478 1898 2482 1902
rect 2486 1898 2490 1902
rect 2486 1838 2490 1842
rect 2486 1808 2490 1812
rect 2470 1788 2474 1792
rect 2454 1768 2458 1772
rect 2454 1738 2458 1742
rect 2462 1708 2466 1712
rect 2486 1728 2490 1732
rect 2478 1618 2482 1622
rect 2398 1518 2402 1522
rect 2390 1508 2394 1512
rect 2422 1508 2426 1512
rect 2414 1448 2418 1452
rect 2390 1428 2394 1432
rect 2422 1428 2426 1432
rect 2382 1418 2386 1422
rect 2406 1378 2410 1382
rect 2382 1338 2386 1342
rect 2374 1298 2378 1302
rect 2374 1288 2378 1292
rect 2398 1308 2402 1312
rect 2382 1268 2386 1272
rect 2366 1078 2370 1082
rect 2406 1298 2410 1302
rect 2398 1238 2402 1242
rect 2454 1538 2458 1542
rect 2478 1468 2482 1472
rect 2446 1448 2450 1452
rect 2454 1448 2458 1452
rect 2470 1388 2474 1392
rect 2478 1378 2482 1382
rect 2462 1368 2466 1372
rect 2470 1318 2474 1322
rect 2430 1268 2434 1272
rect 2438 1268 2442 1272
rect 2438 1258 2442 1262
rect 2430 1198 2434 1202
rect 2538 2003 2542 2007
rect 2545 2003 2546 2007
rect 2546 2003 2549 2007
rect 2566 1978 2570 1982
rect 2538 1803 2542 1807
rect 2545 1803 2546 1807
rect 2546 1803 2549 1807
rect 2510 1798 2514 1802
rect 2558 1798 2562 1802
rect 2550 1778 2554 1782
rect 2518 1748 2522 1752
rect 2550 1688 2554 1692
rect 2558 1678 2562 1682
rect 2518 1658 2522 1662
rect 2534 1658 2538 1662
rect 2526 1628 2530 1632
rect 2574 1818 2578 1822
rect 2622 2438 2626 2442
rect 2670 2328 2674 2332
rect 2646 2298 2650 2302
rect 2662 2238 2666 2242
rect 2638 2018 2642 2022
rect 2590 1818 2594 1822
rect 2538 1603 2542 1607
rect 2545 1603 2546 1607
rect 2546 1603 2549 1607
rect 2590 1748 2594 1752
rect 2606 1748 2610 1752
rect 2614 1718 2618 1722
rect 2614 1678 2618 1682
rect 2590 1648 2594 1652
rect 2526 1598 2530 1602
rect 2582 1598 2586 1602
rect 2510 1578 2514 1582
rect 2598 1628 2602 1632
rect 2502 1558 2506 1562
rect 2558 1538 2562 1542
rect 2534 1528 2538 1532
rect 2558 1528 2562 1532
rect 2502 1398 2506 1402
rect 2486 1218 2490 1222
rect 2486 1168 2490 1172
rect 2478 1158 2482 1162
rect 2478 1148 2482 1152
rect 2406 1138 2410 1142
rect 2438 1088 2442 1092
rect 2414 1078 2418 1082
rect 2430 1078 2434 1082
rect 2430 998 2434 1002
rect 2446 988 2450 992
rect 2478 888 2482 892
rect 2470 878 2474 882
rect 2414 848 2418 852
rect 2414 778 2418 782
rect 2414 688 2418 692
rect 2374 658 2378 662
rect 2334 478 2338 482
rect 2318 268 2322 272
rect 2262 118 2266 122
rect 2286 88 2290 92
rect 2238 58 2242 62
rect 1630 48 1634 52
rect 1798 48 1802 52
rect 2302 178 2306 182
rect 2326 128 2330 132
rect 2334 108 2338 112
rect 2318 98 2322 102
rect 2326 88 2330 92
rect 2334 78 2338 82
rect 2358 348 2362 352
rect 2566 1518 2570 1522
rect 2566 1478 2570 1482
rect 2590 1548 2594 1552
rect 2550 1468 2554 1472
rect 2550 1448 2554 1452
rect 2526 1438 2530 1442
rect 2538 1403 2542 1407
rect 2545 1403 2546 1407
rect 2546 1403 2549 1407
rect 2526 1328 2530 1332
rect 2526 1308 2530 1312
rect 2510 1288 2514 1292
rect 2518 1288 2522 1292
rect 2510 1258 2514 1262
rect 2538 1203 2542 1207
rect 2545 1203 2546 1207
rect 2546 1203 2549 1207
rect 2518 1148 2522 1152
rect 2550 1128 2554 1132
rect 2550 1038 2554 1042
rect 2526 1018 2530 1022
rect 2518 1008 2522 1012
rect 2538 1003 2542 1007
rect 2545 1003 2546 1007
rect 2546 1003 2549 1007
rect 2502 798 2506 802
rect 2462 738 2466 742
rect 2486 728 2490 732
rect 2502 638 2506 642
rect 2470 418 2474 422
rect 2470 378 2474 382
rect 2438 308 2442 312
rect 2462 308 2466 312
rect 2398 268 2402 272
rect 2382 258 2386 262
rect 2538 803 2542 807
rect 2545 803 2546 807
rect 2546 803 2549 807
rect 2526 738 2530 742
rect 2538 603 2542 607
rect 2545 603 2546 607
rect 2546 603 2549 607
rect 2538 403 2542 407
rect 2545 403 2546 407
rect 2546 403 2549 407
rect 2598 1458 2602 1462
rect 2582 1388 2586 1392
rect 2598 1378 2602 1382
rect 2574 1048 2578 1052
rect 2590 1328 2594 1332
rect 2598 1298 2602 1302
rect 2598 1218 2602 1222
rect 2606 1188 2610 1192
rect 2630 1718 2634 1722
rect 2654 2028 2658 2032
rect 2678 2188 2682 2192
rect 2678 1948 2682 1952
rect 2766 2668 2770 2672
rect 2646 1788 2650 1792
rect 2662 1788 2666 1792
rect 2686 1868 2690 1872
rect 2686 1698 2690 1702
rect 2678 1688 2682 1692
rect 2662 1658 2666 1662
rect 2654 1628 2658 1632
rect 2646 1568 2650 1572
rect 2654 1558 2658 1562
rect 2662 1508 2666 1512
rect 2670 1488 2674 1492
rect 2638 1348 2642 1352
rect 2654 1348 2658 1352
rect 2646 1268 2650 1272
rect 2630 1258 2634 1262
rect 2678 1478 2682 1482
rect 2878 2958 2882 2962
rect 2814 2758 2818 2762
rect 2798 2528 2802 2532
rect 2750 2068 2754 2072
rect 2734 2028 2738 2032
rect 2742 1968 2746 1972
rect 2750 1968 2754 1972
rect 2806 2338 2810 2342
rect 2766 1988 2770 1992
rect 2726 1908 2730 1912
rect 2726 1858 2730 1862
rect 2718 1738 2722 1742
rect 2702 1718 2706 1722
rect 2678 1368 2682 1372
rect 2710 1378 2714 1382
rect 2694 1338 2698 1342
rect 2686 1328 2690 1332
rect 2654 1238 2658 1242
rect 2582 978 2586 982
rect 2606 968 2610 972
rect 2574 928 2578 932
rect 2566 908 2570 912
rect 2638 778 2642 782
rect 2630 728 2634 732
rect 2654 1068 2658 1072
rect 2662 938 2666 942
rect 2670 898 2674 902
rect 2758 1848 2762 1852
rect 2734 1708 2738 1712
rect 2758 1678 2762 1682
rect 2742 1578 2746 1582
rect 2750 1558 2754 1562
rect 2750 1528 2754 1532
rect 2734 1518 2738 1522
rect 2726 1508 2730 1512
rect 2702 1248 2706 1252
rect 2758 1478 2762 1482
rect 2742 1448 2746 1452
rect 2750 1418 2754 1422
rect 2742 1368 2746 1372
rect 2742 1328 2746 1332
rect 2734 1298 2738 1302
rect 2742 1258 2746 1262
rect 2774 1568 2778 1572
rect 2758 1308 2762 1312
rect 2710 1148 2714 1152
rect 2718 1128 2722 1132
rect 2742 1118 2746 1122
rect 2758 1108 2762 1112
rect 2798 2038 2802 2042
rect 2822 2578 2826 2582
rect 2854 2538 2858 2542
rect 2838 2478 2842 2482
rect 2822 2278 2826 2282
rect 2814 1978 2818 1982
rect 2798 1758 2802 1762
rect 2814 1638 2818 1642
rect 2870 2578 2874 2582
rect 2886 2728 2890 2732
rect 2934 2938 2938 2942
rect 2942 2588 2946 2592
rect 3042 3103 3046 3107
rect 3049 3103 3050 3107
rect 3050 3103 3053 3107
rect 3502 3278 3506 3282
rect 3302 3268 3306 3272
rect 3510 3268 3514 3272
rect 3118 3258 3122 3262
rect 3094 3248 3098 3252
rect 3102 3158 3106 3162
rect 3042 2903 3046 2907
rect 3049 2903 3050 2907
rect 3050 2903 3053 2907
rect 3126 2888 3130 2892
rect 3150 2868 3154 2872
rect 2918 2498 2922 2502
rect 2862 2248 2866 2252
rect 2870 2028 2874 2032
rect 2894 2318 2898 2322
rect 2958 2478 2962 2482
rect 2918 2108 2922 2112
rect 2902 2058 2906 2062
rect 2862 1988 2866 1992
rect 2870 1978 2874 1982
rect 2854 1898 2858 1902
rect 2846 1878 2850 1882
rect 2846 1858 2850 1862
rect 2830 1718 2834 1722
rect 2838 1548 2842 1552
rect 2798 1528 2802 1532
rect 2798 1438 2802 1442
rect 2766 1078 2770 1082
rect 2678 858 2682 862
rect 2662 708 2666 712
rect 2566 438 2570 442
rect 2502 278 2506 282
rect 2494 268 2498 272
rect 2702 838 2706 842
rect 2710 818 2714 822
rect 2742 828 2746 832
rect 2750 748 2754 752
rect 2662 538 2666 542
rect 2606 468 2610 472
rect 2582 348 2586 352
rect 2558 248 2562 252
rect 2478 238 2482 242
rect 2350 158 2354 162
rect 2366 138 2370 142
rect 2366 108 2370 112
rect 2366 58 2370 62
rect 2486 168 2490 172
rect 2398 138 2402 142
rect 2406 128 2410 132
rect 2406 118 2410 122
rect 2390 68 2394 72
rect 2478 98 2482 102
rect 2538 203 2542 207
rect 2545 203 2546 207
rect 2546 203 2549 207
rect 2526 108 2530 112
rect 2502 88 2506 92
rect 2462 58 2466 62
rect 2686 448 2690 452
rect 2734 478 2738 482
rect 2582 288 2586 292
rect 2694 258 2698 262
rect 2718 228 2722 232
rect 2662 158 2666 162
rect 2582 78 2586 82
rect 2750 148 2754 152
rect 2710 108 2714 112
rect 2750 58 2754 62
rect 2686 38 2690 42
rect 2774 318 2778 322
rect 2774 138 2778 142
rect 2822 1418 2826 1422
rect 2830 1388 2834 1392
rect 2830 1358 2834 1362
rect 2934 2148 2938 2152
rect 2942 2138 2946 2142
rect 2918 1958 2922 1962
rect 2926 1948 2930 1952
rect 2942 1948 2946 1952
rect 3014 2768 3018 2772
rect 3042 2703 3046 2707
rect 3049 2703 3050 2707
rect 3050 2703 3053 2707
rect 3042 2503 3046 2507
rect 3049 2503 3050 2507
rect 3050 2503 3053 2507
rect 2990 2468 2994 2472
rect 3182 2578 3186 2582
rect 3174 2478 3178 2482
rect 3142 2338 3146 2342
rect 2958 2158 2962 2162
rect 2966 2158 2970 2162
rect 3042 2303 3046 2307
rect 3049 2303 3050 2307
rect 3050 2303 3053 2307
rect 3110 2288 3114 2292
rect 3094 2248 3098 2252
rect 2990 2228 2994 2232
rect 2998 2168 3002 2172
rect 3030 2128 3034 2132
rect 3042 2103 3046 2107
rect 3049 2103 3050 2107
rect 3050 2103 3053 2107
rect 3150 2268 3154 2272
rect 3198 2268 3202 2272
rect 3150 2148 3154 2152
rect 3150 2058 3154 2062
rect 3046 2048 3050 2052
rect 3006 2038 3010 2042
rect 2974 1988 2978 1992
rect 3014 1968 3018 1972
rect 3062 1938 3066 1942
rect 2910 1828 2914 1832
rect 2910 1728 2914 1732
rect 2926 1818 2930 1822
rect 2878 1628 2882 1632
rect 2886 1558 2890 1562
rect 2894 1548 2898 1552
rect 2806 1328 2810 1332
rect 2814 1328 2818 1332
rect 2854 1318 2858 1322
rect 2830 1298 2834 1302
rect 2846 1288 2850 1292
rect 2854 1288 2858 1292
rect 2838 1278 2842 1282
rect 2870 1298 2874 1302
rect 2838 1238 2842 1242
rect 2798 538 2802 542
rect 2790 478 2794 482
rect 2790 468 2794 472
rect 2814 1078 2818 1082
rect 2902 1428 2906 1432
rect 2942 1748 2946 1752
rect 2942 1678 2946 1682
rect 2918 1508 2922 1512
rect 2926 1468 2930 1472
rect 2894 1408 2898 1412
rect 2918 1338 2922 1342
rect 2926 1328 2930 1332
rect 2910 1298 2914 1302
rect 2902 1258 2906 1262
rect 2886 1168 2890 1172
rect 2838 688 2842 692
rect 2862 1118 2866 1122
rect 2918 1278 2922 1282
rect 2918 1258 2922 1262
rect 2862 1048 2866 1052
rect 2894 928 2898 932
rect 2862 888 2866 892
rect 2846 548 2850 552
rect 2806 278 2810 282
rect 2798 268 2802 272
rect 2822 258 2826 262
rect 2838 158 2842 162
rect 2830 148 2834 152
rect 2806 128 2810 132
rect 2798 88 2802 92
rect 2902 848 2906 852
rect 2918 1048 2922 1052
rect 2918 968 2922 972
rect 2950 1178 2954 1182
rect 3042 1903 3046 1907
rect 3049 1903 3050 1907
rect 3050 1903 3053 1907
rect 3062 1888 3066 1892
rect 2998 1868 3002 1872
rect 3006 1858 3010 1862
rect 2982 1758 2986 1762
rect 2998 1758 3002 1762
rect 2982 1688 2986 1692
rect 2974 1398 2978 1402
rect 2974 1318 2978 1322
rect 3006 1328 3010 1332
rect 2982 1298 2986 1302
rect 2974 1278 2978 1282
rect 2990 1278 2994 1282
rect 2982 1268 2986 1272
rect 2966 1138 2970 1142
rect 2934 918 2938 922
rect 2926 838 2930 842
rect 2894 658 2898 662
rect 2878 368 2882 372
rect 2982 1148 2986 1152
rect 2950 1008 2954 1012
rect 2966 738 2970 742
rect 2942 348 2946 352
rect 2942 338 2946 342
rect 2870 148 2874 152
rect 2878 128 2882 132
rect 2942 148 2946 152
rect 2934 138 2938 142
rect 2902 118 2906 122
rect 2998 948 3002 952
rect 2974 308 2978 312
rect 3042 1703 3046 1707
rect 3049 1703 3050 1707
rect 3050 1703 3053 1707
rect 3030 1688 3034 1692
rect 3030 1678 3034 1682
rect 3070 1798 3074 1802
rect 3126 1868 3130 1872
rect 3078 1618 3082 1622
rect 3166 1838 3170 1842
rect 3158 1798 3162 1802
rect 3198 2078 3202 2082
rect 3198 1948 3202 1952
rect 3206 1938 3210 1942
rect 3302 3158 3306 3162
rect 3278 2958 3282 2962
rect 3262 2928 3266 2932
rect 3238 2528 3242 2532
rect 3230 2248 3234 2252
rect 3238 2238 3242 2242
rect 3246 2218 3250 2222
rect 3294 2238 3298 2242
rect 3318 3148 3322 3152
rect 3310 2588 3314 2592
rect 3310 2328 3314 2332
rect 3318 2288 3322 2292
rect 3270 1958 3274 1962
rect 3190 1788 3194 1792
rect 3174 1718 3178 1722
rect 3182 1668 3186 1672
rect 3174 1618 3178 1622
rect 3078 1568 3082 1572
rect 3070 1548 3074 1552
rect 3042 1503 3046 1507
rect 3049 1503 3050 1507
rect 3050 1503 3053 1507
rect 3030 1328 3034 1332
rect 3042 1303 3046 1307
rect 3049 1303 3050 1307
rect 3050 1303 3053 1307
rect 3062 1218 3066 1222
rect 3042 1103 3046 1107
rect 3049 1103 3050 1107
rect 3050 1103 3053 1107
rect 3062 928 3066 932
rect 3042 903 3046 907
rect 3049 903 3050 907
rect 3050 903 3053 907
rect 3030 848 3034 852
rect 3086 1378 3090 1382
rect 3110 1268 3114 1272
rect 3086 1258 3090 1262
rect 3166 1608 3170 1612
rect 3158 1588 3162 1592
rect 3102 1138 3106 1142
rect 3102 1008 3106 1012
rect 3086 948 3090 952
rect 3086 878 3090 882
rect 3042 703 3046 707
rect 3049 703 3050 707
rect 3050 703 3053 707
rect 3070 668 3074 672
rect 3070 658 3074 662
rect 3046 638 3050 642
rect 3042 503 3046 507
rect 3049 503 3050 507
rect 3050 503 3053 507
rect 2894 88 2898 92
rect 2950 88 2954 92
rect 2934 68 2938 72
rect 2854 48 2858 52
rect 2974 78 2978 82
rect 2982 48 2986 52
rect 2966 38 2970 42
rect 2974 28 2978 32
rect 3014 148 3018 152
rect 3022 108 3026 112
rect 3070 418 3074 422
rect 3118 848 3122 852
rect 3198 1748 3202 1752
rect 3214 1688 3218 1692
rect 3214 1458 3218 1462
rect 3182 1158 3186 1162
rect 3182 1118 3186 1122
rect 3174 838 3178 842
rect 3166 778 3170 782
rect 3158 688 3162 692
rect 3158 548 3162 552
rect 3182 548 3186 552
rect 3094 478 3098 482
rect 3134 468 3138 472
rect 3110 448 3114 452
rect 3158 368 3162 372
rect 3126 348 3130 352
rect 3134 338 3138 342
rect 3118 328 3122 332
rect 3046 318 3050 322
rect 3042 303 3046 307
rect 3049 303 3050 307
rect 3050 303 3053 307
rect 3046 188 3050 192
rect 3042 103 3046 107
rect 3049 103 3050 107
rect 3050 103 3053 107
rect 3038 68 3042 72
rect 3070 58 3074 62
rect 3030 48 3034 52
rect 3254 1458 3258 1462
rect 3302 2068 3306 2072
rect 3350 2338 3354 2342
rect 3342 2158 3346 2162
rect 3350 2128 3354 2132
rect 3366 3008 3370 3012
rect 3366 2858 3370 2862
rect 3366 2358 3370 2362
rect 3366 2218 3370 2222
rect 3358 2068 3362 2072
rect 3350 2048 3354 2052
rect 3326 1828 3330 1832
rect 3334 1648 3338 1652
rect 3310 1638 3314 1642
rect 3270 1388 3274 1392
rect 3278 1338 3282 1342
rect 3206 948 3210 952
rect 3230 938 3234 942
rect 3230 848 3234 852
rect 3246 668 3250 672
rect 3230 548 3234 552
rect 3206 348 3210 352
rect 3278 1078 3282 1082
rect 3278 938 3282 942
rect 3262 328 3266 332
rect 3110 138 3114 142
rect 3182 128 3186 132
rect 3102 118 3106 122
rect 3102 88 3106 92
rect 3310 1358 3314 1362
rect 3302 1288 3306 1292
rect 3302 1128 3306 1132
rect 3350 1798 3354 1802
rect 3358 1668 3362 1672
rect 3382 2298 3386 2302
rect 3390 1658 3394 1662
rect 3342 1458 3346 1462
rect 3334 1328 3338 1332
rect 3390 1388 3394 1392
rect 3366 1328 3370 1332
rect 3374 1148 3378 1152
rect 3310 1058 3314 1062
rect 3350 1058 3354 1062
rect 3342 1048 3346 1052
rect 3350 968 3354 972
rect 3366 1048 3370 1052
rect 3358 488 3362 492
rect 3334 468 3338 472
rect 3326 448 3330 452
rect 3326 378 3330 382
rect 3318 148 3322 152
rect 3318 68 3322 72
rect 3350 138 3354 142
rect 3390 188 3394 192
rect 3414 2588 3418 2592
rect 3406 2348 3410 2352
rect 3430 2348 3434 2352
rect 3406 1768 3410 1772
rect 3406 1548 3410 1552
rect 3406 1358 3410 1362
rect 3406 1328 3410 1332
rect 3462 3258 3466 3262
rect 3454 3248 3458 3252
rect 3454 2348 3458 2352
rect 3454 2338 3458 2342
rect 3462 2328 3466 2332
rect 3454 2078 3458 2082
rect 3430 1318 3434 1322
rect 3422 958 3426 962
rect 3406 478 3410 482
rect 3478 2358 3482 2362
rect 3486 2168 3490 2172
rect 3470 1638 3474 1642
rect 3446 1548 3450 1552
rect 3478 1338 3482 1342
rect 3478 1278 3482 1282
rect 3502 1908 3506 1912
rect 3534 1908 3538 1912
rect 3518 1698 3522 1702
rect 3510 1658 3514 1662
rect 3510 1578 3514 1582
rect 3462 958 3466 962
rect 3454 588 3458 592
rect 3422 318 3426 322
rect 3366 128 3370 132
rect 3342 78 3346 82
rect 3350 68 3354 72
rect 3470 348 3474 352
rect 3558 2058 3562 2062
rect 3558 1768 3562 1772
rect 3558 1758 3562 1762
rect 3558 1668 3562 1672
rect 3542 1658 3546 1662
rect 3534 1558 3538 1562
rect 3526 1478 3530 1482
rect 3526 1458 3530 1462
rect 3526 998 3530 1002
rect 3486 68 3490 72
rect 3558 1138 3562 1142
rect 2766 8 2770 12
rect 482 3 486 7
rect 489 3 490 7
rect 490 3 493 7
rect 1514 3 1518 7
rect 1521 3 1522 7
rect 1522 3 1525 7
rect 2538 3 2542 7
rect 2545 3 2546 7
rect 2546 3 2549 7
<< metal5 >>
rect 998 3303 1001 3307
rect 997 3302 1002 3303
rect 1007 3302 1008 3307
rect 2030 3303 2033 3307
rect 2029 3302 2034 3303
rect 2039 3302 2040 3307
rect 3046 3303 3049 3307
rect 3045 3302 3050 3303
rect 3055 3302 3056 3307
rect 1138 3298 1142 3301
rect 2170 3288 2238 3291
rect 3502 3282 3505 3287
rect 1538 3268 2182 3271
rect 2186 3268 2310 3271
rect 3306 3268 3510 3271
rect 1426 3258 2030 3261
rect 2770 3258 3118 3261
rect 614 3251 617 3258
rect 3442 3258 3462 3261
rect 614 3248 2214 3251
rect 2514 3248 3094 3251
rect 3454 3242 3457 3248
rect 1506 3238 1846 3241
rect 1054 3232 1057 3238
rect 486 3203 489 3207
rect 485 3202 490 3203
rect 495 3202 496 3207
rect 1518 3203 1521 3207
rect 1517 3202 1522 3203
rect 1527 3202 1528 3207
rect 2542 3203 2545 3207
rect 2541 3202 2546 3203
rect 2551 3202 2552 3207
rect 1106 3188 1878 3191
rect 1658 3168 1710 3171
rect 2498 3158 2702 3161
rect 3106 3158 3302 3161
rect 2786 3148 3318 3151
rect 986 3138 1334 3141
rect 1450 3138 1814 3141
rect 2226 3138 2766 3141
rect 1994 3128 2166 3131
rect 906 3118 1118 3121
rect 2206 3108 2374 3111
rect 998 3103 1001 3107
rect 997 3102 1002 3103
rect 1007 3102 1008 3107
rect 2030 3103 2033 3107
rect 2029 3102 2034 3103
rect 2039 3102 2040 3107
rect 2206 3102 2209 3108
rect 3046 3103 3049 3107
rect 3045 3102 3050 3103
rect 3055 3102 3056 3107
rect 914 3088 1342 3091
rect 2010 3088 2397 3091
rect 946 3078 1118 3081
rect 2106 3068 2182 3071
rect 2442 3068 2502 3071
rect 1726 3062 1729 3068
rect 170 3058 342 3061
rect 578 3058 614 3061
rect 2386 3058 2502 3061
rect 722 3048 1478 3051
rect 1786 3048 1982 3051
rect 1986 3048 2310 3051
rect 338 3038 438 3041
rect 442 3038 1462 3041
rect 1498 3028 1702 3031
rect 1458 3018 2558 3021
rect 3370 3008 3373 3011
rect 486 3003 489 3007
rect 485 3002 490 3003
rect 495 3002 496 3007
rect 1518 3003 1521 3007
rect 1517 3002 1522 3003
rect 1527 3002 1528 3007
rect 2542 3003 2545 3007
rect 2541 3002 2546 3003
rect 2551 3002 2552 3007
rect 1154 2988 1862 2991
rect 2882 2958 3278 2961
rect 818 2948 1182 2951
rect 2058 2948 2182 2951
rect 754 2938 918 2941
rect 994 2938 1062 2941
rect 1482 2938 1814 2941
rect 1826 2938 2022 2941
rect 842 2928 998 2931
rect 1018 2928 1326 2931
rect 1794 2928 1797 2931
rect 1930 2928 2366 2931
rect 2934 2931 2937 2938
rect 2934 2928 3262 2931
rect 234 2918 846 2921
rect 866 2918 974 2921
rect 1618 2918 1654 2921
rect 1770 2918 1821 2921
rect 1866 2918 2086 2921
rect 1130 2908 1622 2911
rect 1626 2908 1878 2911
rect 998 2903 1001 2907
rect 997 2902 1002 2903
rect 1007 2902 1008 2907
rect 2030 2903 2033 2907
rect 2029 2902 2034 2903
rect 2039 2902 2040 2907
rect 3046 2903 3049 2907
rect 3045 2902 3050 2903
rect 3055 2902 3056 2907
rect 938 2888 1294 2891
rect 1850 2888 2078 2891
rect 2394 2888 3126 2891
rect 290 2878 390 2881
rect 554 2878 774 2881
rect 1550 2881 1553 2888
rect 1122 2878 1553 2881
rect 1898 2878 2525 2881
rect 242 2868 510 2871
rect 914 2868 1134 2871
rect 1994 2868 1997 2871
rect 2114 2868 2246 2871
rect 3154 2868 3369 2871
rect 3366 2862 3369 2868
rect 298 2858 374 2861
rect 1658 2858 1846 2861
rect 1946 2858 1990 2861
rect 1994 2858 2206 2861
rect 2482 2858 2558 2861
rect 282 2848 350 2851
rect 1074 2848 1238 2851
rect 1706 2848 1782 2851
rect 1410 2818 2582 2821
rect 486 2803 489 2807
rect 485 2802 490 2803
rect 495 2802 496 2807
rect 1518 2803 1521 2807
rect 1517 2802 1522 2803
rect 1527 2802 1528 2807
rect 1926 2801 1929 2808
rect 2542 2803 2545 2807
rect 2541 2802 2546 2803
rect 2551 2802 2552 2807
rect 1730 2798 1929 2801
rect 386 2788 1566 2791
rect 570 2768 886 2771
rect 890 2768 1366 2771
rect 1802 2768 1870 2771
rect 2378 2768 3014 2771
rect 874 2758 950 2761
rect 2562 2758 2814 2761
rect 186 2748 326 2751
rect 1194 2748 1222 2751
rect 1426 2738 1790 2741
rect 2070 2741 2073 2748
rect 1970 2738 2073 2741
rect 694 2731 697 2738
rect 2866 2738 2889 2741
rect 2886 2732 2889 2738
rect 538 2728 697 2731
rect 1050 2728 1462 2731
rect 2002 2728 2045 2731
rect 2066 2728 2886 2731
rect 450 2718 654 2721
rect 658 2718 742 2721
rect 1330 2718 1438 2721
rect 1450 2718 1582 2721
rect 1730 2718 2126 2721
rect 506 2708 750 2711
rect 1322 2708 2006 2711
rect 998 2703 1001 2707
rect 997 2702 1002 2703
rect 1007 2702 1008 2707
rect 2030 2703 2033 2707
rect 2029 2702 2034 2703
rect 2039 2702 2040 2707
rect 3046 2703 3049 2707
rect 3045 2702 3050 2703
rect 3055 2702 3056 2707
rect 1226 2698 1358 2701
rect 1402 2698 1422 2701
rect 1762 2698 2014 2701
rect 1002 2688 1662 2691
rect 1218 2678 1326 2681
rect 1130 2668 1161 2671
rect 1506 2668 1606 2671
rect 2106 2668 2246 2671
rect 2314 2668 2398 2671
rect 2498 2668 2593 2671
rect 646 2661 649 2668
rect 1158 2662 1161 2668
rect 2590 2662 2593 2668
rect 2766 2662 2769 2668
rect 522 2658 649 2661
rect 778 2658 905 2661
rect 914 2658 942 2661
rect 1210 2658 2366 2661
rect 722 2648 870 2651
rect 902 2651 905 2658
rect 902 2648 1054 2651
rect 1626 2648 2366 2651
rect 2418 2648 2502 2651
rect 394 2638 478 2641
rect 646 2641 649 2648
rect 482 2638 649 2641
rect 850 2638 942 2641
rect 1306 2638 2142 2641
rect 850 2628 1150 2631
rect 1482 2628 1734 2631
rect 2218 2628 2406 2631
rect 1842 2618 2222 2621
rect 1730 2608 1918 2611
rect 2002 2608 2006 2611
rect 486 2603 489 2607
rect 485 2602 490 2603
rect 495 2602 496 2607
rect 1518 2603 1521 2607
rect 1517 2602 1522 2603
rect 1527 2602 1528 2607
rect 2542 2603 2545 2607
rect 2541 2602 2546 2603
rect 2551 2602 2552 2607
rect 1610 2598 2014 2601
rect 442 2588 614 2591
rect 882 2588 926 2591
rect 1402 2588 2406 2591
rect 2514 2588 2942 2591
rect 3314 2588 3414 2591
rect 474 2578 1462 2581
rect 1490 2578 1862 2581
rect 2618 2578 2822 2581
rect 2874 2578 3182 2581
rect 842 2568 974 2571
rect 1138 2568 1150 2571
rect 1154 2568 1622 2571
rect 1698 2568 1774 2571
rect 1898 2568 2134 2571
rect 2430 2571 2433 2578
rect 2202 2568 2433 2571
rect 10 2558 582 2561
rect 778 2558 1078 2561
rect 1086 2561 1089 2568
rect 1086 2558 1214 2561
rect 1218 2558 1606 2561
rect 1618 2558 1766 2561
rect 1786 2558 1902 2561
rect 2206 2552 2209 2558
rect 2590 2552 2593 2558
rect 282 2548 462 2551
rect 618 2548 1118 2551
rect 1130 2548 1133 2551
rect 1258 2548 2190 2551
rect 530 2538 950 2541
rect 1034 2538 1053 2541
rect 1058 2538 1278 2541
rect 1410 2538 2854 2541
rect 202 2528 534 2531
rect 1058 2528 1545 2531
rect 1674 2528 1838 2531
rect 1850 2528 2038 2531
rect 2062 2528 2174 2531
rect 2266 2528 2526 2531
rect 2802 2528 3238 2531
rect 186 2518 374 2521
rect 442 2518 1006 2521
rect 1458 2518 1533 2521
rect 1542 2521 1545 2528
rect 2062 2522 2065 2528
rect 1542 2518 1854 2521
rect 2210 2518 2486 2521
rect 618 2508 942 2511
rect 1226 2508 1638 2511
rect 2442 2508 2461 2511
rect 998 2503 1001 2507
rect 997 2502 1002 2503
rect 1007 2502 1008 2507
rect 2030 2503 2033 2507
rect 2029 2502 2034 2503
rect 2039 2502 2040 2507
rect 3046 2503 3049 2507
rect 3045 2502 3050 2503
rect 3055 2502 3056 2507
rect 1042 2498 1358 2501
rect 1562 2498 1662 2501
rect 2074 2498 2278 2501
rect 2354 2498 2918 2501
rect 218 2488 934 2491
rect 978 2488 1062 2491
rect 1106 2488 2134 2491
rect 474 2478 1262 2481
rect 1442 2478 2838 2481
rect 2962 2478 3174 2481
rect 882 2468 1102 2471
rect 1434 2468 2990 2471
rect 658 2458 830 2461
rect 834 2458 1238 2461
rect 1410 2458 2286 2461
rect 2474 2458 2542 2461
rect 106 2448 598 2451
rect 602 2448 1038 2451
rect 1138 2448 1494 2451
rect 1538 2448 1582 2451
rect 1654 2448 2350 2451
rect 658 2438 1118 2441
rect 1654 2441 1657 2448
rect 1298 2438 1657 2441
rect 1942 2438 2622 2441
rect 418 2428 502 2431
rect 586 2428 798 2431
rect 1942 2431 1945 2438
rect 1370 2428 1945 2431
rect 674 2418 846 2421
rect 890 2418 1390 2421
rect 1410 2418 2526 2421
rect 670 2411 673 2418
rect 506 2408 673 2411
rect 730 2408 822 2411
rect 826 2408 1350 2411
rect 1538 2408 2438 2411
rect 486 2403 489 2407
rect 485 2402 490 2403
rect 495 2402 496 2407
rect 1518 2403 1521 2407
rect 1517 2402 1522 2403
rect 1527 2402 1528 2407
rect 2542 2403 2545 2407
rect 2541 2402 2546 2403
rect 2551 2402 2552 2407
rect 1698 2398 1718 2401
rect 1754 2398 2350 2401
rect 530 2388 966 2391
rect 1026 2388 1270 2391
rect 1490 2388 2310 2391
rect 290 2378 1158 2381
rect 1274 2378 1782 2381
rect 26 2368 574 2371
rect 906 2368 1150 2371
rect 1154 2368 1230 2371
rect 1282 2368 1870 2371
rect 1878 2371 1881 2378
rect 1878 2368 2230 2371
rect 10 2358 622 2361
rect 738 2358 902 2361
rect 1594 2358 1662 2361
rect 1786 2358 1950 2361
rect 1970 2358 2118 2361
rect 3370 2358 3409 2361
rect 394 2348 558 2351
rect 762 2348 958 2351
rect 1010 2348 1478 2351
rect 1658 2348 1742 2351
rect 2334 2351 2337 2358
rect 2106 2348 2337 2351
rect 3406 2352 3409 2358
rect 3474 2358 3478 2361
rect 3434 2348 3454 2351
rect 10 2338 454 2341
rect 578 2338 734 2341
rect 890 2338 1030 2341
rect 1090 2338 1438 2341
rect 1774 2341 1777 2348
rect 1726 2338 1777 2341
rect 2074 2338 2598 2341
rect 2810 2338 3142 2341
rect 3354 2338 3454 2341
rect 542 2332 545 2337
rect 1726 2332 1729 2338
rect 666 2328 782 2331
rect 1194 2328 1709 2331
rect 1754 2328 1830 2331
rect 1946 2328 2270 2331
rect 2498 2328 2502 2331
rect 2674 2328 3310 2331
rect 3458 2328 3462 2331
rect 370 2318 406 2321
rect 410 2318 590 2321
rect 610 2318 1214 2321
rect 1354 2318 1862 2321
rect 1914 2318 1950 2321
rect 1962 2318 2102 2321
rect 2602 2318 2894 2321
rect 722 2308 726 2311
rect 730 2308 798 2311
rect 1250 2308 1294 2311
rect 1898 2308 2006 2311
rect 998 2303 1001 2307
rect 997 2302 1002 2303
rect 1007 2302 1008 2307
rect 2030 2303 2033 2307
rect 2029 2302 2034 2303
rect 2039 2302 2040 2307
rect 3046 2303 3049 2307
rect 3045 2302 3050 2303
rect 3055 2302 3056 2307
rect 1122 2298 1454 2301
rect 2050 2298 2646 2301
rect 3378 2298 3382 2301
rect 986 2288 1286 2291
rect 1522 2288 1830 2291
rect 1834 2288 2102 2291
rect 2170 2288 2270 2291
rect 3114 2288 3318 2291
rect 346 2278 710 2281
rect 730 2278 1014 2281
rect 1062 2278 1414 2281
rect 2026 2278 2142 2281
rect 2170 2278 2574 2281
rect 2598 2278 2822 2281
rect 1062 2272 1065 2278
rect 2598 2272 2601 2278
rect 1258 2268 1430 2271
rect 1530 2268 1582 2271
rect 1722 2268 1725 2271
rect 1730 2268 2094 2271
rect 2114 2268 2198 2271
rect 2202 2268 2382 2271
rect 3154 2268 3198 2271
rect 562 2258 566 2261
rect 1178 2258 1430 2261
rect 2074 2258 2206 2261
rect 14 2248 590 2251
rect 858 2248 1454 2251
rect 2130 2248 2174 2251
rect 2866 2248 3094 2251
rect 3098 2248 3230 2251
rect 14 2242 17 2248
rect 578 2238 670 2241
rect 1130 2238 2662 2241
rect 3242 2238 3294 2241
rect 370 2228 694 2231
rect 1186 2228 1574 2231
rect 2066 2228 2566 2231
rect 546 2218 750 2221
rect 1106 2218 1702 2221
rect 1706 2218 2086 2221
rect 2990 2221 2993 2228
rect 2990 2218 3246 2221
rect 3250 2218 3366 2221
rect 522 2208 1501 2211
rect 1554 2208 1790 2211
rect 2514 2208 2518 2211
rect 486 2203 489 2207
rect 485 2202 490 2203
rect 495 2202 496 2207
rect 1518 2203 1521 2207
rect 1517 2202 1522 2203
rect 1527 2202 1528 2207
rect 2542 2203 2545 2207
rect 2541 2202 2546 2203
rect 2551 2202 2552 2207
rect 682 2198 1070 2201
rect 1658 2198 1846 2201
rect 690 2188 726 2191
rect 858 2188 950 2191
rect 1242 2188 1494 2191
rect 1506 2188 1558 2191
rect 1714 2188 2678 2191
rect 210 2178 1414 2181
rect 1634 2178 1894 2181
rect 2066 2178 2254 2181
rect 1534 2172 1537 2178
rect 586 2168 605 2171
rect 778 2168 1422 2171
rect 1778 2168 2182 2171
rect 2186 2168 2998 2171
rect 3486 2162 3489 2168
rect 554 2158 990 2161
rect 1746 2158 2958 2161
rect 2970 2158 3342 2161
rect 234 2148 582 2151
rect 602 2148 814 2151
rect 930 2148 1841 2151
rect 1850 2148 1958 2151
rect 2938 2148 3150 2151
rect 978 2138 1486 2141
rect 1838 2141 1841 2148
rect 1838 2138 1926 2141
rect 2530 2138 2942 2141
rect 178 2128 717 2131
rect 778 2128 998 2131
rect 1802 2128 2046 2131
rect 3034 2128 3350 2131
rect 1790 2122 1793 2127
rect 1234 2118 1646 2121
rect 1850 2118 2129 2121
rect 2138 2118 2526 2121
rect 650 2108 926 2111
rect 2126 2111 2129 2118
rect 2126 2108 2381 2111
rect 2586 2108 2918 2111
rect 998 2103 1001 2107
rect 997 2102 1002 2103
rect 1007 2102 1008 2107
rect 2030 2103 2033 2107
rect 2029 2102 2034 2103
rect 2039 2102 2040 2107
rect 3046 2103 3049 2107
rect 3045 2102 3050 2103
rect 3055 2102 3056 2107
rect 1386 2098 1758 2101
rect 2058 2098 2134 2101
rect 2206 2092 2209 2097
rect 938 2088 1310 2091
rect 1922 2088 2166 2091
rect 274 2078 526 2081
rect 690 2078 1086 2081
rect 1578 2078 2382 2081
rect 2426 2078 2429 2081
rect 3202 2078 3454 2081
rect 530 2068 598 2071
rect 722 2068 1102 2071
rect 1586 2068 2286 2071
rect 3198 2071 3201 2078
rect 2754 2068 3201 2071
rect 3306 2068 3358 2071
rect 602 2058 798 2061
rect 1410 2058 1726 2061
rect 1738 2058 1741 2061
rect 1906 2058 2062 2061
rect 2178 2058 2182 2061
rect 2906 2058 3150 2061
rect 3154 2058 3558 2061
rect 970 2048 1558 2051
rect 1842 2048 1862 2051
rect 1914 2048 2126 2051
rect 2342 2051 2345 2058
rect 2154 2048 2345 2051
rect 2426 2048 2486 2051
rect 3050 2048 3350 2051
rect 306 2038 878 2041
rect 1474 2038 1582 2041
rect 1594 2038 1702 2041
rect 1770 2038 2294 2041
rect 2802 2038 3006 2041
rect 474 2028 1726 2031
rect 1734 2031 1737 2038
rect 1734 2028 1830 2031
rect 1930 2028 2654 2031
rect 2738 2028 2870 2031
rect 594 2018 606 2021
rect 1026 2018 1038 2021
rect 1106 2018 1310 2021
rect 1506 2018 1654 2021
rect 1682 2018 1773 2021
rect 1786 2018 2638 2021
rect 850 2008 853 2011
rect 1650 2008 1774 2011
rect 1834 2008 1993 2011
rect 486 2003 489 2007
rect 485 2002 490 2003
rect 495 2002 496 2007
rect 1518 2003 1521 2007
rect 1517 2002 1522 2003
rect 1527 2002 1528 2007
rect 658 1998 733 2001
rect 1674 1998 1838 2001
rect 1990 2001 1993 2008
rect 2002 2008 2526 2011
rect 2542 2003 2545 2007
rect 2541 2002 2546 2003
rect 2551 2002 2552 2007
rect 1990 1998 2110 2001
rect 690 1988 1614 1991
rect 1850 1988 2766 1991
rect 2866 1988 2974 1991
rect 82 1978 406 1981
rect 474 1978 534 1981
rect 1042 1978 1949 1981
rect 2202 1978 2566 1981
rect 2818 1978 2870 1981
rect 970 1968 1629 1971
rect 1666 1968 1901 1971
rect 1906 1968 1974 1971
rect 1994 1968 2742 1971
rect 2754 1968 3014 1971
rect 1370 1958 1438 1961
rect 1474 1958 1670 1961
rect 1682 1958 1854 1961
rect 1882 1958 2062 1961
rect 2090 1958 2797 1961
rect 2922 1958 3270 1961
rect 614 1948 942 1951
rect 946 1948 1254 1951
rect 1586 1948 1917 1951
rect 614 1942 617 1948
rect 1922 1948 1942 1951
rect 1954 1948 2077 1951
rect 2098 1948 2102 1951
rect 2306 1948 2309 1951
rect 2682 1948 2926 1951
rect 2946 1948 3198 1951
rect 626 1938 974 1941
rect 1410 1938 1854 1941
rect 2214 1938 2502 1941
rect 3066 1938 3206 1941
rect 954 1928 1086 1931
rect 1554 1928 1646 1931
rect 1654 1928 1718 1931
rect 1726 1928 1782 1931
rect 1786 1928 1789 1931
rect 898 1918 1046 1921
rect 1602 1918 1622 1921
rect 1654 1921 1657 1928
rect 1634 1918 1657 1921
rect 1726 1921 1729 1928
rect 1802 1928 2038 1931
rect 2214 1931 2217 1938
rect 2114 1928 2217 1931
rect 2226 1928 2438 1931
rect 1674 1918 1729 1921
rect 1778 1918 1830 1921
rect 1922 1918 1933 1921
rect 2002 1918 2126 1921
rect 2386 1918 2653 1921
rect 1474 1908 1790 1911
rect 1890 1908 2014 1911
rect 2130 1908 2158 1911
rect 2234 1908 2237 1911
rect 2330 1908 2726 1911
rect 3506 1908 3534 1911
rect 998 1903 1001 1907
rect 997 1902 1002 1903
rect 1007 1902 1008 1907
rect 2030 1903 2033 1907
rect 2029 1902 2034 1903
rect 2039 1902 2040 1907
rect 3046 1903 3049 1907
rect 3045 1902 3050 1903
rect 3055 1902 3056 1907
rect 914 1898 934 1901
rect 1106 1898 1182 1901
rect 1602 1898 1757 1901
rect 1770 1898 1773 1901
rect 1834 1898 1950 1901
rect 2218 1898 2478 1901
rect 2490 1898 2854 1901
rect 194 1888 1265 1891
rect 1274 1888 1769 1891
rect 1778 1888 1894 1891
rect 1898 1888 2222 1891
rect 2242 1888 2253 1891
rect 522 1878 998 1881
rect 1158 1878 1206 1881
rect 1262 1881 1265 1888
rect 1262 1878 1526 1881
rect 1690 1878 1693 1881
rect 1158 1872 1161 1878
rect 1714 1878 1758 1881
rect 1766 1881 1769 1888
rect 2354 1888 3062 1891
rect 1766 1878 2157 1881
rect 2434 1878 2637 1881
rect 2834 1878 2846 1881
rect 2686 1872 2689 1877
rect 562 1868 573 1871
rect 626 1868 637 1871
rect 978 1868 1094 1871
rect 1494 1868 1677 1871
rect 170 1858 398 1861
rect 594 1858 726 1861
rect 1058 1858 1142 1861
rect 1494 1861 1497 1868
rect 1698 1868 1734 1871
rect 1746 1868 1902 1871
rect 1946 1868 2189 1871
rect 2282 1868 2285 1871
rect 3002 1868 3126 1871
rect 1170 1858 1497 1861
rect 1506 1858 1598 1861
rect 1634 1858 1710 1861
rect 1722 1858 1725 1861
rect 1994 1858 2014 1861
rect 2026 1858 2110 1861
rect 2122 1858 2302 1861
rect 2410 1858 2726 1861
rect 2846 1852 2849 1858
rect 3006 1852 3009 1858
rect 458 1848 1374 1851
rect 1506 1848 1654 1851
rect 1706 1848 1750 1851
rect 1858 1848 2278 1851
rect 2286 1848 2758 1851
rect 626 1838 1165 1841
rect 1330 1838 1485 1841
rect 1762 1838 1862 1841
rect 1874 1838 1885 1841
rect 1898 1838 1910 1841
rect 2002 1838 2013 1841
rect 2042 1838 2190 1841
rect 2286 1841 2289 1848
rect 2194 1838 2289 1841
rect 2338 1838 2477 1841
rect 2490 1838 3166 1841
rect 274 1828 654 1831
rect 690 1828 694 1831
rect 754 1828 1078 1831
rect 1082 1828 1118 1831
rect 1122 1828 1334 1831
rect 1346 1828 1349 1831
rect 1474 1828 1997 1831
rect 2026 1828 2061 1831
rect 2074 1828 2153 1831
rect 386 1818 1542 1821
rect 1594 1818 1710 1821
rect 1754 1818 2142 1821
rect 2150 1821 2153 1828
rect 2162 1828 2349 1831
rect 2914 1828 3326 1831
rect 2150 1818 2269 1821
rect 2274 1818 2574 1821
rect 2594 1818 2926 1821
rect 594 1808 909 1811
rect 1074 1808 1462 1811
rect 1538 1808 1686 1811
rect 1778 1808 2061 1811
rect 2090 1808 2486 1811
rect 486 1803 489 1807
rect 485 1802 490 1803
rect 495 1802 496 1807
rect 1518 1803 1521 1807
rect 1517 1802 1522 1803
rect 1527 1802 1528 1807
rect 2542 1803 2545 1807
rect 2541 1802 2546 1803
rect 2551 1802 2552 1807
rect 642 1798 749 1801
rect 962 1798 1502 1801
rect 1618 1798 1833 1801
rect 1842 1798 1934 1801
rect 2002 1798 2230 1801
rect 234 1788 574 1791
rect 1090 1788 1229 1791
rect 1258 1788 1574 1791
rect 1610 1788 1638 1791
rect 1658 1788 1718 1791
rect 1830 1791 1833 1798
rect 2418 1798 2510 1801
rect 2562 1798 3070 1801
rect 3074 1798 3158 1801
rect 3162 1798 3350 1801
rect 1830 1788 2086 1791
rect 2114 1788 2470 1791
rect 2530 1788 2646 1791
rect 2666 1788 3190 1791
rect 434 1778 686 1781
rect 794 1778 1094 1781
rect 1146 1778 1421 1781
rect 1490 1778 1709 1781
rect 1730 1778 1934 1781
rect 1938 1778 2049 1781
rect 2098 1778 2198 1781
rect 2218 1778 2550 1781
rect 458 1768 957 1771
rect 982 1768 990 1771
rect 994 1768 1062 1771
rect 1074 1768 1246 1771
rect 1314 1768 1373 1771
rect 1378 1768 1422 1771
rect 1682 1768 1702 1771
rect 1730 1768 1846 1771
rect 1866 1768 1926 1771
rect 1946 1768 2038 1771
rect 2046 1771 2049 1778
rect 2046 1768 2118 1771
rect 2266 1768 2454 1771
rect 3410 1768 3558 1771
rect 498 1758 1310 1761
rect 1362 1758 1486 1761
rect 1546 1758 1910 1761
rect 1914 1758 2166 1761
rect 2426 1758 2798 1761
rect 3002 1758 3558 1761
rect 290 1748 646 1751
rect 698 1748 1325 1751
rect 138 1738 166 1741
rect 238 1741 241 1748
rect 1378 1748 1437 1751
rect 1506 1748 1790 1751
rect 1794 1748 2086 1751
rect 2138 1748 2518 1751
rect 238 1738 518 1741
rect 650 1738 726 1741
rect 818 1738 1238 1741
rect 1266 1738 1294 1741
rect 1366 1738 1449 1741
rect 2134 1741 2137 1748
rect 2530 1748 2590 1751
rect 2610 1748 2942 1751
rect 2982 1751 2985 1758
rect 2982 1748 3198 1751
rect 1586 1738 2137 1741
rect 466 1728 510 1731
rect 658 1728 870 1731
rect 930 1728 1054 1731
rect 1090 1728 1134 1731
rect 1366 1731 1369 1738
rect 1162 1728 1369 1731
rect 1378 1728 1405 1731
rect 1446 1731 1449 1738
rect 2290 1738 2454 1741
rect 2482 1738 2718 1741
rect 1446 1728 1846 1731
rect 1930 1728 1982 1731
rect 2066 1728 2222 1731
rect 2242 1728 2358 1731
rect 2370 1728 2406 1731
rect 2490 1728 2910 1731
rect 1422 1722 1425 1727
rect 370 1718 590 1721
rect 714 1718 769 1721
rect 858 1718 934 1721
rect 322 1708 542 1711
rect 766 1711 769 1718
rect 962 1718 1198 1721
rect 1210 1718 1382 1721
rect 1434 1718 1518 1721
rect 1602 1718 1798 1721
rect 1818 1718 1821 1721
rect 1954 1718 2109 1721
rect 2122 1718 2398 1721
rect 2434 1718 2609 1721
rect 2618 1718 2621 1721
rect 766 1708 926 1711
rect 1026 1708 1038 1711
rect 1050 1708 1158 1711
rect 1242 1708 1309 1711
rect 1330 1708 2014 1711
rect 2058 1708 2334 1711
rect 2402 1708 2462 1711
rect 2606 1711 2609 1718
rect 2634 1718 2702 1721
rect 2834 1718 3174 1721
rect 2606 1708 2734 1711
rect 998 1703 1001 1707
rect 997 1702 1002 1703
rect 1007 1702 1008 1707
rect 2030 1703 2033 1707
rect 2029 1702 2034 1703
rect 2039 1702 2040 1707
rect 3046 1703 3049 1707
rect 3045 1702 3050 1703
rect 3055 1702 3056 1707
rect 338 1698 557 1701
rect 562 1698 669 1701
rect 714 1698 966 1701
rect 1026 1698 1566 1701
rect 1570 1698 1678 1701
rect 1698 1698 1766 1701
rect 1770 1698 1958 1701
rect 2150 1698 2686 1701
rect 314 1688 766 1691
rect 774 1688 1278 1691
rect 1282 1688 1430 1691
rect 1474 1688 1661 1691
rect 282 1678 621 1681
rect 774 1681 777 1688
rect 1714 1688 1790 1691
rect 1802 1688 1805 1691
rect 2150 1691 2153 1698
rect 3518 1692 3521 1698
rect 1946 1688 2153 1691
rect 2210 1688 2214 1691
rect 2354 1688 2550 1691
rect 2682 1688 2982 1691
rect 3034 1688 3214 1691
rect 682 1678 777 1681
rect 786 1678 1190 1681
rect 1298 1678 1654 1681
rect 1658 1678 1878 1681
rect 1890 1678 1918 1681
rect 1922 1678 2078 1681
rect 2114 1678 2349 1681
rect 2354 1678 2365 1681
rect 2378 1678 2558 1681
rect 2618 1678 2758 1681
rect 2946 1678 3030 1681
rect 866 1668 1038 1671
rect 1066 1668 1118 1671
rect 1170 1668 1449 1671
rect 1458 1668 1510 1671
rect 1562 1668 1581 1671
rect 622 1662 625 1668
rect 402 1658 614 1661
rect 946 1658 974 1661
rect 1058 1658 1166 1661
rect 1186 1658 1277 1661
rect 498 1648 957 1651
rect 970 1648 1125 1651
rect 1294 1651 1297 1658
rect 1314 1658 1389 1661
rect 1410 1658 1438 1661
rect 1446 1661 1449 1668
rect 1594 1668 1757 1671
rect 1770 1668 1789 1671
rect 1826 1668 1837 1671
rect 1858 1668 1958 1671
rect 2066 1668 3182 1671
rect 3362 1668 3558 1671
rect 1446 1658 1982 1661
rect 2002 1658 2518 1661
rect 2538 1658 2662 1661
rect 3514 1658 3542 1661
rect 1138 1648 1297 1651
rect 1306 1648 1718 1651
rect 1730 1648 2046 1651
rect 2050 1648 2190 1651
rect 2274 1648 2590 1651
rect 3390 1651 3393 1658
rect 3338 1648 3393 1651
rect 682 1638 2814 1641
rect 3314 1638 3470 1641
rect 730 1628 774 1631
rect 802 1628 2438 1631
rect 2530 1628 2598 1631
rect 2658 1628 2878 1631
rect 778 1618 1117 1621
rect 1138 1618 1761 1621
rect 1770 1618 2118 1621
rect 2122 1618 2214 1621
rect 2322 1618 2358 1621
rect 2410 1618 2478 1621
rect 3082 1618 3174 1621
rect 666 1608 1398 1611
rect 1410 1608 1478 1611
rect 1554 1608 1557 1611
rect 1714 1608 1725 1611
rect 1758 1611 1761 1618
rect 2366 1612 2369 1618
rect 1758 1608 1790 1611
rect 1794 1608 2334 1611
rect 3170 1608 3501 1611
rect 486 1603 489 1607
rect 485 1602 490 1603
rect 495 1602 496 1607
rect 1518 1603 1521 1607
rect 1517 1602 1522 1603
rect 1527 1602 1528 1607
rect 2542 1603 2545 1607
rect 2541 1602 2546 1603
rect 2551 1602 2552 1607
rect 610 1598 630 1601
rect 882 1598 950 1601
rect 1010 1598 1085 1601
rect 1138 1598 1174 1601
rect 1222 1598 1262 1601
rect 1298 1598 1353 1601
rect 1362 1598 1454 1601
rect 1474 1598 1501 1601
rect 474 1588 1165 1591
rect 1222 1591 1225 1598
rect 1202 1588 1225 1591
rect 1234 1588 1262 1591
rect 1314 1588 1342 1591
rect 338 1578 414 1581
rect 786 1578 1054 1581
rect 1106 1578 1126 1581
rect 1154 1578 1254 1581
rect 1258 1578 1294 1581
rect 1350 1581 1353 1598
rect 1538 1598 1694 1601
rect 1762 1598 1766 1601
rect 1906 1598 2062 1601
rect 2146 1598 2182 1601
rect 2250 1598 2318 1601
rect 2362 1598 2526 1601
rect 2562 1598 2582 1601
rect 1362 1588 1630 1591
rect 1690 1588 1710 1591
rect 1762 1588 1853 1591
rect 1866 1588 1869 1591
rect 1890 1588 1950 1591
rect 1970 1588 1981 1591
rect 1986 1588 2054 1591
rect 2098 1588 3158 1591
rect 1350 1578 1405 1581
rect 1426 1578 1521 1581
rect 1530 1578 1566 1581
rect 1618 1578 1678 1581
rect 1686 1578 1709 1581
rect 594 1568 886 1571
rect 934 1568 1293 1571
rect 474 1558 606 1561
rect 934 1561 937 1568
rect 1394 1568 1414 1571
rect 1442 1568 1510 1571
rect 1518 1571 1521 1578
rect 1686 1572 1689 1578
rect 1754 1578 1870 1581
rect 1938 1578 1958 1581
rect 2018 1578 2105 1581
rect 2114 1578 2150 1581
rect 2154 1578 2326 1581
rect 2338 1578 2422 1581
rect 2514 1578 2742 1581
rect 1518 1568 1582 1571
rect 1714 1568 1966 1571
rect 2010 1568 2061 1571
rect 2102 1571 2105 1578
rect 3490 1578 3510 1581
rect 2102 1568 2150 1571
rect 2166 1568 2353 1571
rect 2362 1568 2477 1571
rect 2166 1562 2169 1568
rect 786 1558 937 1561
rect 946 1558 1149 1561
rect 1170 1558 1286 1561
rect 1322 1558 1574 1561
rect 1658 1558 1734 1561
rect 1778 1558 1853 1561
rect 1890 1558 1990 1561
rect 2010 1558 2013 1561
rect 2050 1558 2118 1561
rect 2138 1558 2166 1561
rect 2210 1558 2302 1561
rect 2350 1561 2353 1568
rect 2486 1568 2646 1571
rect 2778 1568 3078 1571
rect 2486 1561 2489 1568
rect 2350 1558 2489 1561
rect 2506 1558 2654 1561
rect 2754 1558 2886 1561
rect 3362 1558 3534 1561
rect 546 1548 566 1551
rect 1058 1548 1113 1551
rect 286 1538 550 1541
rect 706 1538 717 1541
rect 286 1532 289 1538
rect 962 1538 1030 1541
rect 1110 1541 1113 1548
rect 1122 1548 1142 1551
rect 1186 1548 1309 1551
rect 1330 1548 1334 1551
rect 1378 1548 1437 1551
rect 1458 1548 1494 1551
rect 1506 1548 1590 1551
rect 1602 1548 1625 1551
rect 1634 1548 1766 1551
rect 1810 1548 1862 1551
rect 1110 1538 1213 1541
rect 1234 1538 1342 1541
rect 1378 1538 1422 1541
rect 1458 1538 1478 1541
rect 1498 1538 1613 1541
rect 1622 1541 1625 1548
rect 1922 1548 1934 1551
rect 1978 1548 2070 1551
rect 2082 1548 2278 1551
rect 2290 1548 2573 1551
rect 2594 1548 2765 1551
rect 2842 1548 2894 1551
rect 3074 1548 3406 1551
rect 3450 1548 3469 1551
rect 1622 1538 1886 1541
rect 1898 1538 1982 1541
rect 2058 1538 2222 1541
rect 2306 1538 2454 1541
rect 574 1522 577 1528
rect 594 1528 606 1531
rect 754 1528 1229 1531
rect 1266 1528 2102 1531
rect 2246 1531 2249 1538
rect 2482 1538 2558 1541
rect 2122 1528 2249 1531
rect 2258 1528 2318 1531
rect 2322 1528 2534 1531
rect 2562 1528 2750 1531
rect 2794 1528 2798 1531
rect 162 1518 534 1521
rect 866 1518 886 1521
rect 946 1518 1037 1521
rect 1162 1518 2158 1521
rect 2194 1518 2270 1521
rect 2290 1518 2398 1521
rect 2570 1518 2734 1521
rect 362 1508 365 1511
rect 1066 1508 1101 1511
rect 1234 1508 1329 1511
rect 1338 1508 1374 1511
rect 998 1503 1001 1507
rect 997 1502 1002 1503
rect 1007 1502 1008 1507
rect 1014 1498 1278 1501
rect 1290 1498 1309 1501
rect 1014 1491 1017 1498
rect 1314 1498 1318 1501
rect 1326 1501 1329 1508
rect 1410 1508 1414 1511
rect 1418 1508 1454 1511
rect 1466 1508 2006 1511
rect 2066 1508 2174 1511
rect 2234 1508 2390 1511
rect 2426 1508 2662 1511
rect 2730 1508 2918 1511
rect 2030 1503 2033 1507
rect 2029 1502 2034 1503
rect 2039 1502 2040 1507
rect 3046 1503 3049 1507
rect 3045 1502 3050 1503
rect 3055 1502 3056 1507
rect 1326 1498 1422 1501
rect 1434 1498 1478 1501
rect 1490 1498 1661 1501
rect 1682 1498 1894 1501
rect 1906 1498 1926 1501
rect 1938 1498 2006 1501
rect 2050 1498 2097 1501
rect 2106 1498 2125 1501
rect 138 1488 1017 1491
rect 1122 1488 1182 1491
rect 1218 1488 1606 1491
rect 1634 1488 1878 1491
rect 1890 1488 1949 1491
rect 1994 1488 2077 1491
rect 2094 1491 2097 1498
rect 2162 1498 2206 1501
rect 2250 1498 2285 1501
rect 2306 1498 2334 1501
rect 2354 1498 2358 1501
rect 2094 1488 2321 1491
rect 2346 1488 2493 1491
rect 354 1478 422 1481
rect 450 1478 694 1481
rect 890 1478 893 1481
rect 986 1478 1278 1481
rect 1290 1478 1318 1481
rect 1330 1478 1374 1481
rect 1386 1478 1494 1481
rect 1506 1478 1558 1481
rect 1594 1478 1630 1481
rect 1658 1478 1766 1481
rect 1778 1478 1917 1481
rect 1922 1478 2302 1481
rect 2318 1481 2321 1488
rect 2658 1488 2670 1491
rect 2318 1478 2566 1481
rect 2682 1478 2758 1481
rect 3330 1478 3526 1481
rect 1034 1468 1142 1471
rect 1150 1468 1261 1471
rect 1022 1462 1025 1467
rect 634 1458 998 1461
rect 1150 1461 1153 1468
rect 1282 1468 1329 1471
rect 1338 1468 1614 1471
rect 1034 1458 1153 1461
rect 1194 1458 1206 1461
rect 1218 1458 1246 1461
rect 1250 1458 1270 1461
rect 1326 1461 1329 1468
rect 1634 1468 2013 1471
rect 2042 1468 2045 1471
rect 2122 1468 2262 1471
rect 2354 1468 2478 1471
rect 2554 1468 2926 1471
rect 1326 1458 1389 1461
rect 1426 1458 1518 1461
rect 1546 1458 2302 1461
rect 2322 1458 2598 1461
rect 3218 1458 3254 1461
rect 3346 1458 3526 1461
rect 658 1448 982 1451
rect 1010 1448 1062 1451
rect 1122 1448 1134 1451
rect 1138 1448 1230 1451
rect 1266 1448 1814 1451
rect 1834 1448 1837 1451
rect 1842 1448 2198 1451
rect 2274 1448 2414 1451
rect 2434 1448 2446 1451
rect 2458 1448 2461 1451
rect 2554 1448 2742 1451
rect 402 1438 1390 1441
rect 1394 1438 1422 1441
rect 1474 1438 1478 1441
rect 1538 1438 1606 1441
rect 1618 1438 1654 1441
rect 1658 1438 1709 1441
rect 1738 1438 1757 1441
rect 1778 1438 2214 1441
rect 2386 1438 2526 1441
rect 2578 1438 2798 1441
rect 338 1428 1254 1431
rect 1266 1428 1485 1431
rect 1514 1428 1565 1431
rect 1618 1428 1766 1431
rect 1786 1428 1885 1431
rect 1938 1428 1942 1431
rect 2002 1428 2054 1431
rect 2082 1428 2358 1431
rect 2394 1428 2397 1431
rect 2426 1428 2902 1431
rect 834 1418 845 1421
rect 1002 1418 1046 1421
rect 1058 1418 1094 1421
rect 1202 1418 1421 1421
rect 1506 1418 2030 1421
rect 2034 1418 2078 1421
rect 2114 1418 2134 1421
rect 2138 1418 2382 1421
rect 2422 1418 2750 1421
rect 2754 1418 2822 1421
rect 874 1408 998 1411
rect 1010 1408 1021 1411
rect 1034 1408 1069 1411
rect 1170 1408 1246 1411
rect 1254 1408 1382 1411
rect 1394 1408 1494 1411
rect 1538 1408 1750 1411
rect 1762 1408 1789 1411
rect 486 1403 489 1407
rect 485 1402 490 1403
rect 495 1402 496 1407
rect 746 1398 910 1401
rect 986 1398 1150 1401
rect 1254 1401 1257 1408
rect 1850 1408 2054 1411
rect 2422 1411 2425 1418
rect 2066 1408 2425 1411
rect 2658 1408 2894 1411
rect 1518 1403 1521 1407
rect 1517 1402 1522 1403
rect 1527 1402 1528 1407
rect 2542 1403 2545 1407
rect 2541 1402 2546 1403
rect 2551 1402 2552 1407
rect 1162 1398 1257 1401
rect 1294 1398 1501 1401
rect 1294 1391 1297 1398
rect 1538 1398 1566 1401
rect 1586 1398 1702 1401
rect 1746 1398 1750 1401
rect 1762 1398 1773 1401
rect 1794 1398 1869 1401
rect 1898 1398 2230 1401
rect 2362 1398 2502 1401
rect 2610 1398 2974 1401
rect 450 1388 1297 1391
rect 1306 1388 1341 1391
rect 1354 1388 1870 1391
rect 1874 1388 2365 1391
rect 2474 1388 2573 1391
rect 2586 1388 2830 1391
rect 3274 1388 3390 1391
rect 354 1378 1062 1381
rect 1066 1378 1462 1381
rect 1506 1378 1894 1381
rect 1970 1378 2086 1381
rect 2226 1378 2406 1381
rect 2434 1378 2478 1381
rect 2602 1378 2621 1381
rect 2714 1378 3086 1381
rect 858 1368 893 1371
rect 954 1368 1086 1371
rect 1098 1368 1214 1371
rect 1234 1368 1325 1371
rect 1378 1368 1558 1371
rect 1562 1368 1822 1371
rect 1838 1368 1846 1371
rect 218 1358 230 1361
rect 514 1358 518 1361
rect 594 1358 1325 1361
rect 1342 1361 1345 1368
rect 1342 1358 1366 1361
rect 1490 1358 1598 1361
rect 1618 1358 1677 1361
rect 1838 1361 1841 1368
rect 1874 1368 1990 1371
rect 2106 1368 2230 1371
rect 2242 1368 2366 1371
rect 2466 1368 2678 1371
rect 2706 1368 2742 1371
rect 1698 1358 1841 1361
rect 1850 1358 1870 1361
rect 1898 1358 1942 1361
rect 2018 1358 2222 1361
rect 2242 1358 2270 1361
rect 2282 1358 2350 1361
rect 2370 1358 2830 1361
rect 3314 1358 3406 1361
rect 1438 1352 1441 1357
rect 650 1348 966 1351
rect 978 1348 982 1351
rect 1050 1348 1270 1351
rect 1298 1348 1358 1351
rect 1370 1348 1389 1351
rect 530 1338 957 1341
rect 1022 1341 1025 1348
rect 1526 1348 1581 1351
rect 970 1338 1025 1341
rect 1034 1338 1101 1341
rect 1154 1338 1206 1341
rect 1234 1338 1310 1341
rect 1330 1338 1382 1341
rect 1526 1341 1529 1348
rect 1590 1348 1597 1351
rect 1402 1338 1529 1341
rect 1590 1341 1593 1348
rect 1714 1348 1822 1351
rect 1882 1348 1926 1351
rect 1938 1348 1949 1351
rect 1954 1348 1997 1351
rect 2034 1348 2078 1351
rect 2090 1348 2173 1351
rect 2238 1351 2241 1357
rect 2186 1348 2241 1351
rect 2266 1348 2638 1351
rect 1694 1342 1697 1347
rect 1586 1338 1593 1341
rect 1602 1338 1606 1341
rect 1666 1338 1678 1341
rect 1770 1338 1806 1341
rect 1890 1338 1981 1341
rect 2242 1338 2365 1341
rect 2386 1338 2525 1341
rect 2654 1341 2657 1348
rect 2578 1338 2657 1341
rect 2698 1338 2809 1341
rect 2922 1338 3278 1341
rect 3482 1338 3485 1341
rect 2094 1332 2097 1337
rect 2742 1332 2745 1338
rect 2806 1332 2809 1338
rect 370 1328 830 1331
rect 914 1328 942 1331
rect 978 1328 1390 1331
rect 1506 1328 1686 1331
rect 1690 1328 1750 1331
rect 1770 1328 1878 1331
rect 1890 1328 2006 1331
rect 2018 1328 2046 1331
rect 2114 1328 2182 1331
rect 2306 1328 2526 1331
rect 2594 1328 2686 1331
rect 2818 1328 2926 1331
rect 3002 1328 3006 1331
rect 3034 1328 3334 1331
rect 3370 1328 3406 1331
rect 730 1318 966 1321
rect 978 1318 990 1321
rect 1010 1318 1037 1321
rect 1122 1318 1158 1321
rect 1306 1318 1709 1321
rect 1070 1312 1073 1318
rect 1722 1318 1725 1321
rect 1778 1318 1862 1321
rect 1882 1318 1902 1321
rect 1982 1312 1985 1318
rect 2018 1318 2094 1321
rect 2274 1318 2285 1321
rect 2474 1318 2854 1321
rect 2978 1318 3430 1321
rect 418 1308 670 1311
rect 858 1308 974 1311
rect 1026 1308 1038 1311
rect 1154 1308 1501 1311
rect 1510 1308 1734 1311
rect 1754 1308 1942 1311
rect 998 1303 1001 1307
rect 997 1302 1002 1303
rect 1007 1302 1008 1307
rect 1510 1301 1513 1308
rect 2058 1308 2061 1311
rect 2030 1303 2033 1307
rect 2029 1302 2034 1303
rect 2039 1302 2040 1307
rect 2046 1302 2049 1308
rect 2122 1308 2237 1311
rect 2250 1308 2398 1311
rect 2530 1308 2758 1311
rect 3046 1303 3049 1307
rect 3045 1302 3050 1303
rect 3055 1302 3056 1307
rect 1042 1298 1513 1301
rect 1546 1298 1702 1301
rect 1722 1298 1782 1301
rect 1826 1298 1918 1301
rect 858 1288 1478 1291
rect 1490 1288 1550 1291
rect 1570 1288 1629 1291
rect 1666 1288 1758 1291
rect 1798 1291 1801 1298
rect 1970 1298 1974 1301
rect 2106 1298 2166 1301
rect 2178 1298 2374 1301
rect 2410 1298 2413 1301
rect 2578 1298 2598 1301
rect 2738 1298 2749 1301
rect 2834 1298 2870 1301
rect 2914 1298 2982 1301
rect 1798 1288 1902 1291
rect 1946 1288 2077 1291
rect 2098 1288 2158 1291
rect 2210 1288 2289 1291
rect 2378 1288 2510 1291
rect 2522 1288 2846 1291
rect 2858 1288 3302 1291
rect 2286 1282 2289 1288
rect 618 1278 782 1281
rect 786 1278 870 1281
rect 962 1278 1110 1281
rect 1138 1278 1238 1281
rect 626 1268 742 1271
rect 786 1268 862 1271
rect 946 1268 1021 1271
rect 1034 1268 1206 1271
rect 1242 1268 1262 1271
rect 1310 1271 1313 1278
rect 1410 1278 1705 1281
rect 1786 1278 2182 1281
rect 1298 1268 1313 1271
rect 658 1258 801 1261
rect 850 1258 950 1261
rect 970 1258 1053 1261
rect 798 1252 801 1258
rect 1090 1258 1278 1261
rect 1298 1258 1309 1261
rect 1342 1261 1345 1268
rect 1426 1268 1470 1271
rect 1546 1268 1638 1271
rect 1642 1268 1677 1271
rect 1702 1271 1705 1278
rect 2306 1278 2350 1281
rect 2362 1278 2838 1281
rect 2922 1278 2974 1281
rect 2994 1278 3478 1281
rect 1702 1268 2150 1271
rect 2154 1268 2382 1271
rect 2418 1268 2430 1271
rect 2442 1268 2445 1271
rect 2642 1268 2646 1271
rect 2986 1268 3110 1271
rect 2510 1262 2513 1267
rect 1330 1258 1345 1261
rect 1362 1258 1422 1261
rect 1434 1258 1437 1261
rect 1542 1258 1902 1261
rect 1954 1258 2054 1261
rect 2098 1258 2262 1261
rect 2290 1258 2438 1261
rect 210 1248 246 1251
rect 306 1248 398 1251
rect 458 1248 686 1251
rect 1002 1248 1022 1251
rect 1042 1248 1085 1251
rect 1542 1251 1545 1258
rect 2594 1258 2630 1261
rect 2746 1258 2902 1261
rect 2922 1258 3086 1261
rect 1098 1248 1545 1251
rect 1554 1248 2118 1251
rect 2146 1248 2157 1251
rect 2242 1248 2702 1251
rect 450 1238 1102 1241
rect 1114 1238 1197 1241
rect 1210 1238 1422 1241
rect 1450 1238 2230 1241
rect 2306 1238 2317 1241
rect 2402 1238 2654 1241
rect 2834 1238 2838 1241
rect 234 1228 846 1231
rect 862 1228 1246 1231
rect 1250 1228 1597 1231
rect 862 1221 865 1228
rect 1626 1228 1670 1231
rect 1698 1228 1702 1231
rect 1714 1228 1741 1231
rect 1786 1228 2206 1231
rect 2338 1228 2573 1231
rect 466 1218 865 1221
rect 874 1218 1838 1221
rect 1874 1218 1974 1221
rect 1986 1218 2038 1221
rect 2082 1218 2350 1221
rect 2362 1218 2486 1221
rect 2602 1218 3062 1221
rect 730 1208 926 1211
rect 946 1208 949 1211
rect 978 1208 990 1211
rect 1026 1208 1494 1211
rect 1554 1208 1590 1211
rect 1698 1208 1830 1211
rect 1842 1208 2190 1211
rect 2626 1208 2685 1211
rect 486 1203 489 1207
rect 485 1202 490 1203
rect 495 1202 496 1207
rect 1518 1203 1521 1207
rect 1517 1202 1522 1203
rect 1527 1202 1528 1207
rect 1646 1202 1649 1207
rect 2542 1203 2545 1207
rect 2541 1202 2546 1203
rect 2551 1202 2552 1207
rect 754 1198 941 1201
rect 966 1198 1502 1201
rect 966 1191 969 1198
rect 1538 1198 1566 1201
rect 1730 1198 1758 1201
rect 1762 1198 2070 1201
rect 2082 1198 2430 1201
rect 390 1188 969 1191
rect 978 1188 1118 1191
rect 1194 1188 1262 1191
rect 1266 1188 1325 1191
rect 390 1182 393 1188
rect 1338 1188 1389 1191
rect 1394 1188 1430 1191
rect 1458 1188 1742 1191
rect 1754 1188 1894 1191
rect 1898 1188 2606 1191
rect 834 1178 1046 1181
rect 1106 1178 1229 1181
rect 1242 1178 1245 1181
rect 1290 1178 1814 1181
rect 1954 1178 2093 1181
rect 2178 1178 2950 1181
rect 578 1168 846 1171
rect 954 1168 1094 1171
rect 1122 1168 1318 1171
rect 1330 1168 1341 1171
rect 1386 1168 1438 1171
rect 1490 1168 1542 1171
rect 1586 1168 1769 1171
rect 1778 1168 1966 1171
rect 2010 1168 2182 1171
rect 2274 1168 2429 1171
rect 462 1162 465 1167
rect 690 1158 1022 1161
rect 1066 1158 1222 1161
rect 1242 1158 1277 1161
rect 1306 1158 1325 1161
rect 1410 1158 1702 1161
rect 1714 1158 1734 1161
rect 1746 1158 1757 1161
rect 1766 1161 1769 1168
rect 2490 1168 2886 1171
rect 1766 1158 2137 1161
rect 2146 1158 2478 1161
rect 402 1148 510 1151
rect 714 1148 749 1151
rect 826 1148 838 1151
rect 914 1148 1037 1151
rect 1074 1148 1133 1151
rect 1154 1148 1225 1151
rect 1250 1148 1342 1151
rect 1346 1148 1373 1151
rect 1222 1142 1225 1148
rect 1466 1148 1581 1151
rect 1602 1148 1869 1151
rect 1938 1148 1965 1151
rect 1986 1148 2062 1151
rect 2074 1148 2109 1151
rect 2134 1151 2137 1158
rect 2134 1148 2237 1151
rect 2482 1148 2518 1151
rect 2522 1148 2710 1151
rect 3182 1151 3185 1158
rect 2986 1148 3185 1151
rect 3378 1148 3561 1151
rect 3558 1142 3561 1148
rect 930 1138 1086 1141
rect 1114 1138 1181 1141
rect 670 1132 673 1138
rect 1258 1138 1277 1141
rect 1306 1138 1309 1141
rect 1338 1138 1366 1141
rect 1378 1138 1382 1141
rect 1394 1138 1542 1141
rect 1578 1138 1622 1141
rect 1650 1138 1798 1141
rect 1818 1138 2174 1141
rect 2178 1138 2294 1141
rect 2410 1138 2605 1141
rect 2970 1138 3102 1141
rect 842 1128 861 1131
rect 874 1128 1126 1131
rect 1138 1128 1281 1131
rect 730 1118 1126 1121
rect 1146 1118 1174 1121
rect 1186 1118 1206 1121
rect 1278 1121 1281 1128
rect 1318 1128 1486 1131
rect 1318 1121 1321 1128
rect 1570 1128 1597 1131
rect 1618 1128 1665 1131
rect 1690 1128 1790 1131
rect 1810 1128 1878 1131
rect 1890 1128 1958 1131
rect 1662 1122 1665 1128
rect 2066 1128 2078 1131
rect 2234 1128 2350 1131
rect 2554 1128 2557 1131
rect 2722 1128 3302 1131
rect 1278 1118 1321 1121
rect 1330 1118 1421 1121
rect 1474 1118 1645 1121
rect 666 1108 982 1111
rect 1034 1108 1134 1111
rect 1254 1111 1257 1118
rect 1682 1118 1709 1121
rect 1722 1118 1990 1121
rect 2014 1118 2310 1121
rect 2354 1118 2742 1121
rect 2866 1118 3182 1121
rect 1146 1108 1257 1111
rect 1266 1108 1294 1111
rect 1322 1108 1325 1111
rect 1346 1108 1453 1111
rect 1458 1108 1598 1111
rect 1650 1108 1670 1111
rect 1682 1108 1806 1111
rect 1834 1108 1873 1111
rect 1882 1108 1934 1111
rect 998 1103 1001 1107
rect 997 1102 1002 1103
rect 1007 1102 1008 1107
rect 714 1098 814 1101
rect 818 1098 925 1101
rect 1042 1098 1190 1101
rect 1202 1098 1702 1101
rect 1714 1098 1846 1101
rect 1870 1101 1873 1108
rect 1954 1108 1958 1111
rect 2014 1111 2017 1118
rect 1970 1108 2017 1111
rect 2066 1108 2077 1111
rect 2090 1108 2758 1111
rect 2030 1103 2033 1107
rect 2029 1102 2034 1103
rect 2039 1102 2040 1107
rect 3046 1103 3049 1107
rect 3045 1102 3050 1103
rect 3055 1102 3056 1107
rect 1870 1098 2006 1101
rect 2050 1098 2413 1101
rect 626 1088 870 1091
rect 970 1088 1062 1091
rect 1114 1088 1149 1091
rect 1162 1088 1341 1091
rect 1354 1088 1405 1091
rect 1442 1088 1478 1091
rect 1490 1088 1622 1091
rect 1698 1088 1773 1091
rect 1778 1088 1806 1091
rect 1818 1088 2166 1091
rect 2178 1088 2254 1091
rect 2290 1088 2294 1091
rect 2442 1088 2653 1091
rect 786 1078 1030 1081
rect 1042 1078 1165 1081
rect 1170 1078 1270 1081
rect 1298 1078 1334 1081
rect 1346 1078 1374 1081
rect 1458 1078 1558 1081
rect 1602 1078 1718 1081
rect 1722 1078 1837 1081
rect 1898 1078 2126 1081
rect 2250 1078 2350 1081
rect 2370 1078 2397 1081
rect 2434 1078 2766 1081
rect 2818 1078 3278 1081
rect 618 1068 910 1071
rect 962 1068 1142 1071
rect 1154 1068 1334 1071
rect 1370 1068 1462 1071
rect 1474 1068 1485 1071
rect 1618 1068 1670 1071
rect 1674 1068 1734 1071
rect 1746 1068 1805 1071
rect 1810 1068 2013 1071
rect 2414 1071 2417 1078
rect 2210 1068 2417 1071
rect 2658 1068 2861 1071
rect 234 1058 1022 1061
rect 622 1052 625 1058
rect 1162 1058 1438 1061
rect 1442 1058 1822 1061
rect 1858 1058 1910 1061
rect 1930 1058 2134 1061
rect 2162 1058 2349 1061
rect 3314 1058 3350 1061
rect 1118 1052 1121 1057
rect 442 1048 582 1051
rect 658 1048 838 1051
rect 850 1048 877 1051
rect 978 1048 982 1051
rect 1130 1048 1213 1051
rect 1234 1048 1526 1051
rect 1538 1048 2070 1051
rect 2098 1048 2574 1051
rect 2866 1048 2918 1051
rect 3346 1048 3366 1051
rect 506 1038 718 1041
rect 738 1038 1286 1041
rect 1322 1038 1462 1041
rect 1474 1038 1613 1041
rect 1618 1038 1630 1041
rect 1650 1038 1741 1041
rect 1754 1038 1902 1041
rect 1938 1038 1958 1041
rect 1986 1038 2174 1041
rect 2194 1038 2550 1041
rect 674 1028 733 1031
rect 746 1028 877 1031
rect 882 1028 2022 1031
rect 2066 1028 2109 1031
rect 2114 1028 2205 1031
rect 2226 1028 2326 1031
rect 914 1018 974 1021
rect 1010 1018 1245 1021
rect 1258 1018 1277 1021
rect 1282 1018 1318 1021
rect 1346 1018 1670 1021
rect 1690 1018 2526 1021
rect 798 1012 801 1017
rect 946 1008 1174 1011
rect 1202 1008 1246 1011
rect 1274 1008 1414 1011
rect 1498 1008 1502 1011
rect 1594 1008 1694 1011
rect 486 1003 489 1007
rect 485 1002 490 1003
rect 495 1002 496 1007
rect 1518 1003 1521 1007
rect 1517 1002 1522 1003
rect 1527 1002 1528 1007
rect 1582 1002 1585 1008
rect 1746 1008 2518 1011
rect 2954 1008 3102 1011
rect 2542 1003 2545 1007
rect 2541 1002 2546 1003
rect 2551 1002 2552 1007
rect 834 998 846 1001
rect 914 998 1069 1001
rect 1210 998 1502 1001
rect 1666 998 1981 1001
rect 2050 998 2262 1001
rect 2274 998 2430 1001
rect 610 988 1182 991
rect 1218 988 1222 991
rect 1234 988 1257 991
rect 10 978 502 981
rect 962 978 1245 981
rect 1254 981 1257 988
rect 1266 988 1277 991
rect 1330 988 1422 991
rect 1442 988 1693 991
rect 1698 988 2446 991
rect 3526 991 3529 998
rect 3522 988 3529 991
rect 1254 978 1469 981
rect 1490 978 1862 981
rect 1906 978 1933 981
rect 1954 978 1998 981
rect 2018 978 2278 981
rect 2290 978 2582 981
rect 402 968 822 971
rect 826 968 862 971
rect 874 968 1022 971
rect 1130 968 1254 971
rect 1282 968 1550 971
rect 1634 968 2606 971
rect 2922 968 3350 971
rect 394 958 470 961
rect 842 958 982 961
rect 1114 958 1406 961
rect 1046 951 1049 958
rect 1474 958 1590 961
rect 1602 958 1645 961
rect 1682 958 1838 961
rect 1850 958 2022 961
rect 2050 958 2118 961
rect 2130 958 2174 961
rect 2210 958 2230 961
rect 3426 958 3462 961
rect 658 948 1049 951
rect 1058 948 1193 951
rect 1202 948 1726 951
rect 1738 948 1757 951
rect 626 938 957 941
rect 978 938 1062 941
rect 1082 938 1182 941
rect 1190 941 1193 948
rect 1930 948 1958 951
rect 1978 948 2062 951
rect 2354 948 2998 951
rect 3090 948 3206 951
rect 1190 938 1246 941
rect 1298 938 1302 941
rect 1314 938 1469 941
rect 1490 938 1886 941
rect 1938 938 1942 941
rect 1954 938 2302 941
rect 2666 938 2685 941
rect 3234 938 3278 941
rect 466 928 1206 931
rect 1330 928 1406 931
rect 1506 928 1789 931
rect 1834 928 2214 931
rect 2450 928 2574 931
rect 2898 928 3062 931
rect 706 918 710 921
rect 786 918 1214 921
rect 1266 918 1294 921
rect 1338 918 1357 921
rect 1370 918 1494 921
rect 1550 918 1558 921
rect 1562 918 1702 921
rect 1714 918 1718 921
rect 1882 918 1966 921
rect 2018 918 2934 921
rect 866 908 982 911
rect 862 901 865 908
rect 1026 908 1142 911
rect 1154 908 1262 911
rect 1298 908 1302 911
rect 1346 908 1614 911
rect 1674 908 1677 911
rect 1746 908 2013 911
rect 2074 908 2077 911
rect 2098 908 2566 911
rect 998 903 1001 907
rect 997 902 1002 903
rect 1007 902 1008 907
rect 2030 903 2033 907
rect 2029 902 2034 903
rect 2039 902 2040 907
rect 3046 903 3049 907
rect 3045 902 3050 903
rect 3055 902 3056 907
rect 746 898 865 901
rect 1042 898 1206 901
rect 1218 898 1302 901
rect 1322 898 1405 901
rect 1474 898 1750 901
rect 1802 898 1913 901
rect 578 888 638 891
rect 802 888 1166 891
rect 1250 888 1390 891
rect 1426 888 1565 891
rect 1586 888 1725 891
rect 1730 888 1798 891
rect 1910 891 1913 898
rect 1922 898 1950 901
rect 2050 898 2086 901
rect 2162 898 2670 901
rect 1910 888 2014 891
rect 2102 891 2105 898
rect 2026 888 2105 891
rect 2178 888 2478 891
rect 2850 888 2862 891
rect 722 878 1046 881
rect 1050 878 1118 881
rect 1186 878 1198 881
rect 1234 878 1289 881
rect 1298 878 1702 881
rect 1730 878 1937 881
rect 1946 878 2206 881
rect 2474 878 3086 881
rect 802 868 813 871
rect 946 868 966 871
rect 1002 868 1245 871
rect 122 858 342 861
rect 870 861 873 868
rect 1286 871 1289 878
rect 1286 868 1485 871
rect 1506 868 1926 871
rect 1934 871 1937 878
rect 1934 868 1966 871
rect 2074 868 2238 871
rect 2266 868 2310 871
rect 870 858 877 861
rect 962 858 1053 861
rect 1114 858 1206 861
rect 1218 858 1478 861
rect 1490 858 1857 861
rect 1866 858 2086 861
rect 2682 858 2905 861
rect 466 848 558 851
rect 762 848 838 851
rect 930 848 1374 851
rect 1402 848 1429 851
rect 1442 848 1638 851
rect 1650 848 1782 851
rect 1834 848 1846 851
rect 1854 851 1857 858
rect 2902 852 2905 858
rect 1854 848 1934 851
rect 2042 848 2414 851
rect 2906 848 3030 851
rect 3122 848 3230 851
rect 178 838 286 841
rect 714 838 717 841
rect 866 838 2702 841
rect 2930 838 3174 841
rect 594 828 953 831
rect 354 818 622 821
rect 950 821 953 828
rect 1094 828 1142 831
rect 1154 828 1278 831
rect 1094 821 1097 828
rect 1314 828 1318 831
rect 1354 828 1510 831
rect 1514 828 1918 831
rect 1994 828 2742 831
rect 950 818 1097 821
rect 1170 818 1206 821
rect 1218 818 1326 821
rect 1330 818 1870 821
rect 1914 818 2030 821
rect 2050 818 2710 821
rect 666 808 809 811
rect 818 808 1286 811
rect 1290 808 1406 811
rect 486 803 489 807
rect 485 802 490 803
rect 495 802 496 807
rect 786 798 797 801
rect 806 801 809 808
rect 1570 808 2150 811
rect 2186 808 2206 811
rect 1518 803 1521 807
rect 1517 802 1522 803
rect 1527 802 1528 807
rect 2542 803 2545 807
rect 2541 802 2546 803
rect 2551 802 2552 807
rect 806 798 1181 801
rect 1210 798 1502 801
rect 1562 798 1686 801
rect 1698 798 1758 801
rect 1794 798 2093 801
rect 2146 798 2502 801
rect 546 788 654 791
rect 770 788 1158 791
rect 1170 788 1238 791
rect 1250 788 1513 791
rect 1522 788 2062 791
rect 2066 788 2182 791
rect 738 778 966 781
rect 970 778 1478 781
rect 1510 781 1513 788
rect 1510 778 1670 781
rect 1690 778 1766 781
rect 1906 778 2414 781
rect 2642 778 3166 781
rect 458 768 1182 771
rect 1258 768 1337 771
rect 1346 768 2062 771
rect 2122 768 2230 771
rect 2338 768 2701 771
rect 314 758 606 761
rect 978 758 990 761
rect 1186 758 1309 761
rect 1334 761 1337 768
rect 1334 758 1389 761
rect 1394 758 1462 761
rect 1490 758 1990 761
rect 2002 758 2142 761
rect 2750 752 2753 757
rect 786 748 790 751
rect 1162 748 1342 751
rect 1354 748 1598 751
rect 1722 748 1725 751
rect 546 738 830 741
rect 842 738 1117 741
rect 1138 738 1318 741
rect 1338 738 1430 741
rect 1734 741 1737 748
rect 1746 748 1846 751
rect 1938 748 2278 751
rect 1546 738 1737 741
rect 1858 738 1950 741
rect 1970 738 2014 741
rect 2058 738 2158 741
rect 2282 738 2462 741
rect 2530 738 2966 741
rect 282 728 878 731
rect 882 728 909 731
rect 930 728 1246 731
rect 1282 728 1286 731
rect 1306 728 1406 731
rect 1498 728 1997 731
rect 2018 728 2198 731
rect 2202 728 2301 731
rect 2490 728 2630 731
rect 362 718 606 721
rect 610 718 669 721
rect 882 718 1222 721
rect 1226 718 2294 721
rect 250 708 638 711
rect 642 708 718 711
rect 770 708 974 711
rect 1082 708 1254 711
rect 1266 708 1470 711
rect 1490 708 1790 711
rect 2074 708 2662 711
rect 998 703 1001 707
rect 997 702 1002 703
rect 1007 702 1008 707
rect 2030 703 2033 707
rect 2029 702 2034 703
rect 2039 702 2040 707
rect 3046 703 3049 707
rect 3045 702 3050 703
rect 3055 702 3056 707
rect 314 698 365 701
rect 370 698 718 701
rect 890 698 893 701
rect 1074 698 1142 701
rect 1186 698 1390 701
rect 1410 698 1518 701
rect 1522 698 1533 701
rect 1586 698 1614 701
rect 1698 698 1782 701
rect 338 688 678 691
rect 714 688 1134 691
rect 1170 688 1501 691
rect 1530 688 1574 691
rect 1578 688 1709 691
rect 1714 688 1822 691
rect 1870 691 1873 698
rect 1870 688 2414 691
rect 2842 688 3158 691
rect 602 678 950 681
rect 986 678 1078 681
rect 1090 678 1245 681
rect 1282 678 1501 681
rect 1514 678 1782 681
rect 1818 678 2045 681
rect 2090 678 2173 681
rect 274 668 509 671
rect 514 668 910 671
rect 1130 668 1286 671
rect 1338 668 1341 671
rect 1458 668 1502 671
rect 1770 668 2150 671
rect 3074 668 3246 671
rect 130 658 590 661
rect 834 658 910 661
rect 1026 658 1277 661
rect 1298 658 1438 661
rect 1490 658 1693 661
rect 1714 658 1790 661
rect 1826 658 1933 661
rect 2074 658 2374 661
rect 2898 658 3070 661
rect 718 652 721 657
rect 306 648 598 651
rect 890 648 1182 651
rect 1202 648 1241 651
rect 386 638 454 641
rect 786 638 934 641
rect 978 638 1038 641
rect 1058 638 1214 641
rect 1238 641 1241 648
rect 1250 648 1485 651
rect 1506 648 1702 651
rect 1738 648 1854 651
rect 2002 648 2078 651
rect 1238 638 1325 641
rect 1934 641 1937 648
rect 1422 638 1937 641
rect 2506 638 3046 641
rect 606 632 609 637
rect 754 628 1101 631
rect 1202 628 1270 631
rect 1406 631 1409 638
rect 1314 628 1409 631
rect 1422 632 1425 638
rect 1474 628 2254 631
rect 202 618 422 621
rect 570 618 685 621
rect 882 618 1166 621
rect 1178 618 1190 621
rect 1194 618 1486 621
rect 1850 618 1878 621
rect 1922 618 2302 621
rect 1550 612 1553 617
rect 866 608 1037 611
rect 1114 608 1310 611
rect 1322 608 1502 611
rect 1954 608 2166 611
rect 486 603 489 607
rect 485 602 490 603
rect 495 602 496 607
rect 1518 603 1521 607
rect 1517 602 1522 603
rect 1527 602 1528 607
rect 2542 603 2545 607
rect 2541 602 2546 603
rect 2551 602 2552 607
rect 674 598 926 601
rect 930 598 1030 601
rect 1106 598 1278 601
rect 1282 598 1486 601
rect 1898 598 2086 601
rect 514 588 790 591
rect 802 588 877 591
rect 898 588 1086 591
rect 1106 588 3454 591
rect 798 582 801 587
rect 938 578 1006 581
rect 1050 578 1110 581
rect 1138 578 1390 581
rect 910 571 913 578
rect 1410 578 1661 581
rect 910 568 1318 571
rect 1338 568 1622 571
rect 506 558 742 561
rect 818 558 937 561
rect 970 558 1133 561
rect 934 552 937 558
rect 1146 558 1294 561
rect 1314 558 1425 561
rect 1818 558 1821 561
rect 1422 552 1425 558
rect 402 548 550 551
rect 554 548 734 551
rect 842 548 925 551
rect 978 548 1102 551
rect 1122 548 1166 551
rect 1186 548 1302 551
rect 1314 548 1405 551
rect 2850 548 3158 551
rect 3186 548 3230 551
rect 242 538 470 541
rect 826 538 1142 541
rect 1178 538 1278 541
rect 1330 538 1406 541
rect 1970 538 2221 541
rect 2666 538 2798 541
rect 290 528 854 531
rect 1298 528 1718 531
rect 442 518 878 521
rect 1098 518 1334 521
rect 1378 518 1390 521
rect 1410 518 2141 521
rect 250 508 942 511
rect 1026 508 1798 511
rect 1938 508 1949 511
rect 998 503 1001 507
rect 997 502 1002 503
rect 1007 502 1008 507
rect 2030 503 2033 507
rect 2029 502 2034 503
rect 2039 502 2040 507
rect 3046 503 3049 507
rect 3045 502 3050 503
rect 3055 502 3056 507
rect 522 498 973 501
rect 1026 498 1830 501
rect 410 488 766 491
rect 778 488 1414 491
rect 1426 488 3358 491
rect 458 478 686 481
rect 714 478 1494 481
rect 1746 478 2174 481
rect 2226 478 2334 481
rect 2738 478 2790 481
rect 3098 478 3406 481
rect 634 468 1341 471
rect 1346 468 1454 471
rect 2610 468 2790 471
rect 3138 468 3334 471
rect 818 458 1422 461
rect 1570 458 1774 461
rect 2686 452 2689 457
rect 370 448 950 451
rect 3114 448 3326 451
rect 610 438 1006 441
rect 1138 438 1654 441
rect 1922 438 2006 441
rect 2010 438 2566 441
rect 890 428 1254 431
rect 1266 428 1590 431
rect 1618 428 1918 431
rect 626 418 1021 421
rect 1042 418 2077 421
rect 2474 418 3070 421
rect 850 408 1230 411
rect 486 403 489 407
rect 485 402 490 403
rect 495 402 496 407
rect 1518 403 1521 407
rect 1517 402 1522 403
rect 1527 402 1528 407
rect 2542 403 2545 407
rect 2541 402 2546 403
rect 2551 402 2552 407
rect 618 398 1438 401
rect 754 388 1862 391
rect 482 378 774 381
rect 1170 378 1270 381
rect 1274 378 2470 381
rect 3330 378 3437 381
rect 594 368 1958 371
rect 2882 368 3158 371
rect 594 358 654 361
rect 914 358 934 361
rect 962 358 1158 361
rect 1214 351 1217 358
rect 1146 348 1217 351
rect 1706 348 1774 351
rect 1778 348 1838 351
rect 2362 348 2582 351
rect 2946 348 3126 351
rect 3210 348 3470 351
rect 590 342 593 347
rect 546 338 582 341
rect 2946 338 3134 341
rect 474 328 542 331
rect 546 328 621 331
rect 642 328 662 331
rect 674 328 1110 331
rect 2010 328 2118 331
rect 3122 328 3262 331
rect 394 318 454 321
rect 458 318 1030 321
rect 2018 318 2214 321
rect 2770 318 2774 321
rect 3050 318 3422 321
rect 802 308 846 311
rect 1026 308 1422 311
rect 1842 308 1942 311
rect 2162 308 2438 311
rect 2466 308 2974 311
rect 998 303 1001 307
rect 997 302 1002 303
rect 1007 302 1008 307
rect 2030 303 2033 307
rect 2029 302 2034 303
rect 2039 302 2040 307
rect 3046 303 3049 307
rect 3045 302 3050 303
rect 3055 302 3056 307
rect 1330 288 1478 291
rect 1482 288 1806 291
rect 1834 288 2582 291
rect 930 278 1110 281
rect 1114 278 1430 281
rect 1474 278 1598 281
rect 1682 278 1814 281
rect 1866 278 2502 281
rect 2506 278 2806 281
rect 1702 272 1705 278
rect 114 268 278 271
rect 1314 268 1686 271
rect 1762 268 1806 271
rect 1978 268 2062 271
rect 2066 268 2134 271
rect 2322 268 2398 271
rect 2498 268 2798 271
rect 634 258 1022 261
rect 1106 258 1142 261
rect 1578 258 1766 261
rect 2090 258 2238 261
rect 2386 258 2621 261
rect 2698 258 2822 261
rect 810 248 2558 251
rect 610 238 1126 241
rect 1186 238 1310 241
rect 1826 238 1982 241
rect 2170 238 2478 241
rect 690 228 926 231
rect 1274 228 2718 231
rect 698 218 886 221
rect 890 218 1222 221
rect 626 208 934 211
rect 486 203 489 207
rect 485 202 490 203
rect 495 202 496 207
rect 1518 203 1521 207
rect 1517 202 1522 203
rect 1527 202 1528 207
rect 2542 203 2545 207
rect 2541 202 2546 203
rect 2551 202 2552 207
rect 698 188 701 191
rect 882 188 1254 191
rect 3050 188 3390 191
rect 706 178 718 181
rect 954 178 1174 181
rect 1986 178 2302 181
rect 202 168 742 171
rect 778 168 833 171
rect 842 168 926 171
rect 986 168 1134 171
rect 1138 168 2486 171
rect 830 162 833 168
rect 562 158 801 161
rect 850 158 1334 161
rect 2066 158 2094 161
rect 2122 158 2185 161
rect 2354 158 2662 161
rect 2666 158 2838 161
rect 546 148 662 151
rect 798 151 801 158
rect 2182 152 2185 158
rect 798 148 1390 151
rect 1394 148 1438 151
rect 1802 148 2142 151
rect 2754 148 2830 151
rect 2874 148 2942 151
rect 3018 148 3318 151
rect 130 138 726 141
rect 770 138 1318 141
rect 1810 138 2366 141
rect 2402 138 2774 141
rect 2938 138 3110 141
rect 738 128 1502 131
rect 1802 128 2326 131
rect 2410 128 2806 131
rect 2870 128 2878 131
rect 2882 128 3182 131
rect 3350 131 3353 138
rect 3350 128 3366 131
rect 442 118 942 121
rect 1106 118 2262 121
rect 2410 118 2902 121
rect 2906 118 3102 121
rect 378 108 446 111
rect 566 108 670 111
rect 1026 108 1342 111
rect 1482 108 1710 111
rect 2146 108 2334 111
rect 2370 108 2526 111
rect 2714 108 3022 111
rect 566 102 569 108
rect 998 103 1001 107
rect 997 102 1002 103
rect 1007 102 1008 107
rect 2030 103 2033 107
rect 2029 102 2034 103
rect 2039 102 2040 107
rect 3046 103 3049 107
rect 3045 102 3050 103
rect 3055 102 3056 107
rect 370 98 566 101
rect 626 98 814 101
rect 818 98 825 101
rect 1306 98 1374 101
rect 1890 98 2014 101
rect 2322 98 2478 101
rect 354 88 686 91
rect 706 88 1246 91
rect 1290 88 1350 91
rect 1434 88 2286 91
rect 2330 88 2502 91
rect 2802 88 2894 91
rect 2954 88 3102 91
rect 114 78 605 81
rect 610 78 758 81
rect 786 78 838 81
rect 842 78 926 81
rect 1186 78 1494 81
rect 1802 78 1918 81
rect 1978 78 2062 81
rect 2338 78 2582 81
rect 2978 78 3342 81
rect 3486 72 3489 77
rect 434 68 870 71
rect 1098 68 2006 71
rect 2226 68 2390 71
rect 2938 68 3038 71
rect 3322 68 3325 71
rect 3354 68 3357 71
rect 562 58 721 61
rect 1010 58 1142 61
rect 1234 58 1350 61
rect 1354 58 1438 61
rect 1626 58 2238 61
rect 2370 58 2462 61
rect 2754 58 3070 61
rect 490 48 710 51
rect 718 51 721 58
rect 718 48 1038 51
rect 1222 48 1230 51
rect 1234 48 1470 51
rect 1634 48 1798 51
rect 2858 48 2982 51
rect 2986 48 3030 51
rect 706 38 790 41
rect 2690 38 2966 41
rect 730 28 1110 31
rect 1114 28 2974 31
rect 650 18 1014 21
rect 2766 12 2769 17
rect 486 3 489 7
rect 485 2 490 3
rect 495 2 496 7
rect 1518 3 1521 7
rect 1517 2 1522 3
rect 1527 2 1528 7
rect 2542 3 2545 7
rect 2541 2 2546 3
rect 2551 2 2552 7
<< m6contact >>
rect 992 3303 994 3307
rect 994 3303 997 3307
rect 1002 3303 1005 3307
rect 1005 3303 1007 3307
rect 992 3302 997 3303
rect 1002 3302 1007 3303
rect 2024 3303 2026 3307
rect 2026 3303 2029 3307
rect 2034 3303 2037 3307
rect 2037 3303 2039 3307
rect 2024 3302 2029 3303
rect 2034 3302 2039 3303
rect 3040 3303 3042 3307
rect 3042 3303 3045 3307
rect 3050 3303 3053 3307
rect 3053 3303 3055 3307
rect 3040 3302 3045 3303
rect 3050 3302 3055 3303
rect 1133 3297 1138 3302
rect 3501 3287 3506 3292
rect 3437 3257 3442 3262
rect 3453 3237 3458 3242
rect 1053 3227 1058 3232
rect 480 3203 482 3207
rect 482 3203 485 3207
rect 490 3203 493 3207
rect 493 3203 495 3207
rect 480 3202 485 3203
rect 490 3202 495 3203
rect 1512 3203 1514 3207
rect 1514 3203 1517 3207
rect 1522 3203 1525 3207
rect 1525 3203 1527 3207
rect 1512 3202 1517 3203
rect 1522 3202 1527 3203
rect 2536 3203 2538 3207
rect 2538 3203 2541 3207
rect 2546 3203 2549 3207
rect 2549 3203 2551 3207
rect 2536 3202 2541 3203
rect 2546 3202 2551 3203
rect 992 3103 994 3107
rect 994 3103 997 3107
rect 1002 3103 1005 3107
rect 1005 3103 1007 3107
rect 992 3102 997 3103
rect 1002 3102 1007 3103
rect 2024 3103 2026 3107
rect 2026 3103 2029 3107
rect 2034 3103 2037 3107
rect 2037 3103 2039 3107
rect 2024 3102 2029 3103
rect 2034 3102 2039 3103
rect 3040 3103 3042 3107
rect 3042 3103 3045 3107
rect 3050 3103 3053 3107
rect 3053 3103 3055 3107
rect 3040 3102 3045 3103
rect 3050 3102 3055 3103
rect 2397 3087 2402 3092
rect 1725 3057 1730 3062
rect 3373 3007 3378 3012
rect 480 3003 482 3007
rect 482 3003 485 3007
rect 490 3003 493 3007
rect 493 3003 495 3007
rect 480 3002 485 3003
rect 490 3002 495 3003
rect 1512 3003 1514 3007
rect 1514 3003 1517 3007
rect 1522 3003 1525 3007
rect 1525 3003 1527 3007
rect 1512 3002 1517 3003
rect 1522 3002 1527 3003
rect 2536 3003 2538 3007
rect 2538 3003 2541 3007
rect 2546 3003 2549 3007
rect 2549 3003 2551 3007
rect 2536 3002 2541 3003
rect 2546 3002 2551 3003
rect 1821 2937 1826 2942
rect 1797 2927 1802 2932
rect 1821 2917 1826 2922
rect 992 2903 994 2907
rect 994 2903 997 2907
rect 1002 2903 1005 2907
rect 1005 2903 1007 2907
rect 992 2902 997 2903
rect 1002 2902 1007 2903
rect 2024 2903 2026 2907
rect 2026 2903 2029 2907
rect 2034 2903 2037 2907
rect 2037 2903 2039 2907
rect 2024 2902 2029 2903
rect 2034 2902 2039 2903
rect 3040 2903 3042 2907
rect 3042 2903 3045 2907
rect 3050 2903 3053 2907
rect 3053 2903 3055 2907
rect 3040 2902 3045 2903
rect 3050 2902 3055 2903
rect 2525 2877 2530 2882
rect 1997 2867 2002 2872
rect 480 2803 482 2807
rect 482 2803 485 2807
rect 490 2803 493 2807
rect 493 2803 495 2807
rect 480 2802 485 2803
rect 490 2802 495 2803
rect 1512 2803 1514 2807
rect 1514 2803 1517 2807
rect 1522 2803 1525 2807
rect 1525 2803 1527 2807
rect 1512 2802 1517 2803
rect 1522 2802 1527 2803
rect 2536 2803 2538 2807
rect 2538 2803 2541 2807
rect 2546 2803 2549 2807
rect 2549 2803 2551 2807
rect 2536 2802 2541 2803
rect 2546 2802 2551 2803
rect 2861 2737 2866 2742
rect 2045 2727 2050 2732
rect 992 2703 994 2707
rect 994 2703 997 2707
rect 1002 2703 1005 2707
rect 1005 2703 1007 2707
rect 992 2702 997 2703
rect 1002 2702 1007 2703
rect 2024 2703 2026 2707
rect 2026 2703 2029 2707
rect 2034 2703 2037 2707
rect 2037 2703 2039 2707
rect 2024 2702 2029 2703
rect 2034 2702 2039 2703
rect 3040 2703 3042 2707
rect 3042 2703 3045 2707
rect 3050 2703 3053 2707
rect 3053 2703 3055 2707
rect 3040 2702 3045 2703
rect 3050 2702 3055 2703
rect 2765 2657 2770 2662
rect 1997 2607 2002 2612
rect 480 2603 482 2607
rect 482 2603 485 2607
rect 490 2603 493 2607
rect 493 2603 495 2607
rect 480 2602 485 2603
rect 490 2602 495 2603
rect 1512 2603 1514 2607
rect 1514 2603 1517 2607
rect 1522 2603 1525 2607
rect 1525 2603 1527 2607
rect 1512 2602 1517 2603
rect 1522 2602 1527 2603
rect 2536 2603 2538 2607
rect 2538 2603 2541 2607
rect 2546 2603 2549 2607
rect 2549 2603 2551 2607
rect 2536 2602 2541 2603
rect 2546 2602 2551 2603
rect 1133 2547 1138 2552
rect 2205 2547 2210 2552
rect 2589 2547 2594 2552
rect 1053 2537 1058 2542
rect 1533 2517 1538 2522
rect 2461 2507 2466 2512
rect 992 2503 994 2507
rect 994 2503 997 2507
rect 1002 2503 1005 2507
rect 1005 2503 1007 2507
rect 992 2502 997 2503
rect 1002 2502 1007 2503
rect 2024 2503 2026 2507
rect 2026 2503 2029 2507
rect 2034 2503 2037 2507
rect 2037 2503 2039 2507
rect 2024 2502 2029 2503
rect 2034 2502 2039 2503
rect 3040 2503 3042 2507
rect 3042 2503 3045 2507
rect 3050 2503 3053 2507
rect 3053 2503 3055 2507
rect 3040 2502 3045 2503
rect 3050 2502 3055 2503
rect 1533 2407 1538 2412
rect 480 2403 482 2407
rect 482 2403 485 2407
rect 490 2403 493 2407
rect 493 2403 495 2407
rect 480 2402 485 2403
rect 490 2402 495 2403
rect 1512 2403 1514 2407
rect 1514 2403 1517 2407
rect 1522 2403 1525 2407
rect 1525 2403 1527 2407
rect 1512 2402 1517 2403
rect 1522 2402 1527 2403
rect 2536 2403 2538 2407
rect 2538 2403 2541 2407
rect 2546 2403 2549 2407
rect 2549 2403 2551 2407
rect 2536 2402 2541 2403
rect 2546 2402 2551 2403
rect 3469 2357 3474 2362
rect 541 2337 546 2342
rect 1709 2327 1714 2332
rect 2493 2327 2498 2332
rect 3453 2327 3458 2332
rect 717 2307 722 2312
rect 992 2303 994 2307
rect 994 2303 997 2307
rect 1002 2303 1005 2307
rect 1005 2303 1007 2307
rect 992 2302 997 2303
rect 1002 2302 1007 2303
rect 2024 2303 2026 2307
rect 2026 2303 2029 2307
rect 2034 2303 2037 2307
rect 2037 2303 2039 2307
rect 2024 2302 2029 2303
rect 2034 2302 2039 2303
rect 3040 2303 3042 2307
rect 3042 2303 3045 2307
rect 3050 2303 3053 2307
rect 3053 2303 3055 2307
rect 3040 2302 3045 2303
rect 3050 2302 3055 2303
rect 3373 2297 3378 2302
rect 1725 2267 1730 2272
rect 557 2257 562 2262
rect 2061 2227 2066 2232
rect 541 2217 546 2222
rect 1501 2207 1506 2212
rect 2509 2207 2514 2212
rect 480 2203 482 2207
rect 482 2203 485 2207
rect 490 2203 493 2207
rect 493 2203 495 2207
rect 480 2202 485 2203
rect 490 2202 495 2203
rect 1512 2203 1514 2207
rect 1514 2203 1517 2207
rect 1522 2203 1525 2207
rect 1525 2203 1527 2207
rect 1512 2202 1517 2203
rect 1522 2202 1527 2203
rect 2536 2203 2538 2207
rect 2538 2203 2541 2207
rect 2546 2203 2549 2207
rect 2549 2203 2551 2207
rect 2536 2202 2541 2203
rect 2546 2202 2551 2203
rect 1501 2187 1506 2192
rect 1709 2187 1714 2192
rect 605 2167 610 2172
rect 1533 2167 1538 2172
rect 3485 2157 3490 2162
rect 717 2127 722 2132
rect 1789 2127 1794 2132
rect 2381 2107 2386 2112
rect 992 2103 994 2107
rect 994 2103 997 2107
rect 1002 2103 1005 2107
rect 1005 2103 1007 2107
rect 992 2102 997 2103
rect 1002 2102 1007 2103
rect 2024 2103 2026 2107
rect 2026 2103 2029 2107
rect 2034 2103 2037 2107
rect 2037 2103 2039 2107
rect 2024 2102 2029 2103
rect 2034 2102 2039 2103
rect 3040 2103 3042 2107
rect 3042 2103 3045 2107
rect 3050 2103 3053 2107
rect 3053 2103 3055 2107
rect 3040 2102 3045 2103
rect 3050 2102 3055 2103
rect 2205 2097 2210 2102
rect 2429 2077 2434 2082
rect 1581 2067 1586 2072
rect 1405 2057 1410 2062
rect 1741 2057 1746 2062
rect 2173 2057 2178 2062
rect 1837 2047 1842 2052
rect 589 2017 594 2022
rect 1677 2017 1682 2022
rect 1773 2017 1778 2022
rect 853 2007 858 2012
rect 1645 2007 1650 2012
rect 480 2003 482 2007
rect 482 2003 485 2007
rect 490 2003 493 2007
rect 493 2003 495 2007
rect 480 2002 485 2003
rect 490 2002 495 2003
rect 1512 2003 1514 2007
rect 1514 2003 1517 2007
rect 1522 2003 1525 2007
rect 1525 2003 1527 2007
rect 1512 2002 1517 2003
rect 1522 2002 1527 2003
rect 733 1997 738 2002
rect 1997 2007 2002 2012
rect 2536 2003 2538 2007
rect 2538 2003 2541 2007
rect 2546 2003 2549 2007
rect 2549 2003 2551 2007
rect 2536 2002 2541 2003
rect 2546 2002 2551 2003
rect 1037 1977 1042 1982
rect 1949 1977 1954 1982
rect 1629 1967 1634 1972
rect 1661 1967 1666 1972
rect 1901 1967 1906 1972
rect 2797 1957 2802 1962
rect 1917 1947 1922 1952
rect 1949 1947 1954 1952
rect 2077 1947 2082 1952
rect 2093 1947 2098 1952
rect 2309 1947 2314 1952
rect 893 1917 898 1922
rect 1597 1917 1602 1922
rect 1789 1927 1794 1932
rect 2221 1927 2226 1932
rect 1773 1917 1778 1922
rect 1933 1917 1938 1922
rect 2653 1917 2658 1922
rect 2125 1907 2130 1912
rect 2237 1907 2242 1912
rect 992 1903 994 1907
rect 994 1903 997 1907
rect 1002 1903 1005 1907
rect 1005 1903 1007 1907
rect 992 1902 997 1903
rect 1002 1902 1007 1903
rect 2024 1903 2026 1907
rect 2026 1903 2029 1907
rect 2034 1903 2037 1907
rect 2037 1903 2039 1907
rect 2024 1902 2029 1903
rect 2034 1902 2039 1903
rect 3040 1903 3042 1907
rect 3042 1903 3045 1907
rect 3050 1903 3053 1907
rect 3053 1903 3055 1907
rect 3040 1902 3045 1903
rect 3050 1902 3055 1903
rect 909 1897 914 1902
rect 1101 1897 1106 1902
rect 1757 1897 1762 1902
rect 1773 1897 1778 1902
rect 1693 1877 1698 1882
rect 1709 1877 1714 1882
rect 2253 1887 2258 1892
rect 2349 1887 2354 1892
rect 2157 1877 2162 1882
rect 2637 1877 2642 1882
rect 2685 1877 2690 1882
rect 2829 1877 2834 1882
rect 573 1867 578 1872
rect 637 1867 642 1872
rect 973 1867 978 1872
rect 1053 1857 1058 1862
rect 1165 1857 1170 1862
rect 1677 1867 1682 1872
rect 2189 1867 2194 1872
rect 2285 1867 2290 1872
rect 1725 1857 1730 1862
rect 1501 1847 1506 1852
rect 621 1837 626 1842
rect 1165 1837 1170 1842
rect 1485 1837 1490 1842
rect 1757 1838 1758 1842
rect 1758 1838 1762 1842
rect 1757 1837 1762 1838
rect 1885 1837 1890 1842
rect 2013 1837 2018 1842
rect 2845 1847 2850 1852
rect 3005 1847 3010 1852
rect 2477 1837 2482 1842
rect 685 1827 690 1832
rect 749 1827 754 1832
rect 1349 1827 1354 1832
rect 1469 1827 1474 1832
rect 1997 1827 2002 1832
rect 2061 1827 2066 1832
rect 2157 1827 2162 1832
rect 2349 1827 2354 1832
rect 2269 1817 2274 1822
rect 909 1807 914 1812
rect 1069 1807 1074 1812
rect 2061 1807 2066 1812
rect 480 1803 482 1807
rect 482 1803 485 1807
rect 490 1803 493 1807
rect 493 1803 495 1807
rect 480 1802 485 1803
rect 490 1802 495 1803
rect 1512 1803 1514 1807
rect 1514 1803 1517 1807
rect 1522 1803 1525 1807
rect 1525 1803 1527 1807
rect 1512 1802 1517 1803
rect 1522 1802 1527 1803
rect 2536 1803 2538 1807
rect 2538 1803 2541 1807
rect 2546 1803 2549 1807
rect 2549 1803 2551 1807
rect 2536 1802 2541 1803
rect 2546 1802 2551 1803
rect 749 1797 754 1802
rect 957 1797 962 1802
rect 1229 1787 1234 1792
rect 2413 1797 2418 1802
rect 2109 1787 2114 1792
rect 2525 1787 2530 1792
rect 1421 1777 1426 1782
rect 1485 1777 1490 1782
rect 1709 1777 1714 1782
rect 1725 1777 1730 1782
rect 957 1767 962 1772
rect 1373 1767 1378 1772
rect 1677 1767 1682 1772
rect 1725 1767 1730 1772
rect 1325 1747 1330 1752
rect 1437 1747 1442 1752
rect 1261 1737 1266 1742
rect 2525 1747 2530 1752
rect 461 1727 466 1732
rect 925 1727 930 1732
rect 1085 1727 1090 1732
rect 1405 1727 1410 1732
rect 1421 1727 1426 1732
rect 2285 1737 2290 1742
rect 2477 1737 2482 1742
rect 2365 1727 2370 1732
rect 957 1717 962 1722
rect 1821 1717 1826 1722
rect 1949 1717 1954 1722
rect 2109 1717 2114 1722
rect 1309 1707 1314 1712
rect 2397 1707 2402 1712
rect 2621 1717 2626 1722
rect 992 1703 994 1707
rect 994 1703 997 1707
rect 1002 1703 1005 1707
rect 1005 1703 1007 1707
rect 992 1702 997 1703
rect 1002 1702 1007 1703
rect 2024 1703 2026 1707
rect 2026 1703 2029 1707
rect 2034 1703 2037 1707
rect 2037 1703 2039 1707
rect 2024 1702 2029 1703
rect 2034 1702 2039 1703
rect 3040 1703 3042 1707
rect 3042 1703 3045 1707
rect 3050 1703 3053 1707
rect 3053 1703 3055 1707
rect 3040 1702 3045 1703
rect 3050 1702 3055 1703
rect 557 1697 562 1702
rect 669 1697 674 1702
rect 1021 1697 1026 1702
rect 1661 1688 1662 1692
rect 1662 1688 1666 1692
rect 621 1677 626 1682
rect 1661 1687 1666 1688
rect 1709 1687 1714 1692
rect 1805 1687 1810 1692
rect 2205 1687 2210 1692
rect 3517 1687 3522 1692
rect 2349 1677 2354 1682
rect 2365 1677 2370 1682
rect 621 1657 626 1662
rect 941 1657 946 1662
rect 1181 1657 1186 1662
rect 1277 1657 1282 1662
rect 957 1647 962 1652
rect 1125 1647 1130 1652
rect 1309 1657 1314 1662
rect 1389 1657 1394 1662
rect 1581 1667 1586 1672
rect 1757 1667 1762 1672
rect 1789 1667 1794 1672
rect 1837 1667 1842 1672
rect 1853 1667 1858 1672
rect 2061 1667 2066 1672
rect 1997 1657 2002 1662
rect 1301 1647 1306 1652
rect 797 1627 802 1632
rect 1117 1617 1122 1622
rect 1557 1607 1562 1612
rect 1725 1607 1730 1612
rect 2365 1607 2370 1612
rect 3501 1607 3506 1612
rect 480 1603 482 1607
rect 482 1603 485 1607
rect 490 1603 493 1607
rect 493 1603 495 1607
rect 480 1602 485 1603
rect 490 1602 495 1603
rect 1512 1603 1514 1607
rect 1514 1603 1517 1607
rect 1522 1603 1525 1607
rect 1525 1603 1527 1607
rect 1512 1602 1517 1603
rect 1522 1602 1527 1603
rect 2536 1603 2538 1607
rect 2538 1603 2541 1607
rect 2546 1603 2549 1607
rect 2549 1603 2551 1607
rect 2536 1602 2541 1603
rect 2546 1602 2551 1603
rect 605 1597 610 1602
rect 877 1597 882 1602
rect 1085 1597 1090 1602
rect 1165 1587 1170 1592
rect 1229 1587 1234 1592
rect 1309 1587 1314 1592
rect 1149 1577 1154 1582
rect 1501 1597 1506 1602
rect 1757 1597 1762 1602
rect 2141 1597 2146 1602
rect 2557 1597 2562 1602
rect 1757 1587 1762 1592
rect 1853 1587 1858 1592
rect 1869 1587 1874 1592
rect 1885 1587 1890 1592
rect 1981 1587 1986 1592
rect 1405 1577 1410 1582
rect 1421 1577 1426 1582
rect 1293 1567 1298 1572
rect 1389 1567 1394 1572
rect 1437 1567 1442 1572
rect 1709 1577 1714 1582
rect 1933 1577 1938 1582
rect 2061 1567 2066 1572
rect 3485 1577 3490 1582
rect 1149 1557 1154 1562
rect 1853 1557 1858 1562
rect 2013 1557 2018 1562
rect 2477 1567 2482 1572
rect 3357 1557 3362 1562
rect 717 1537 722 1542
rect 1117 1547 1122 1552
rect 1181 1547 1186 1552
rect 1309 1547 1314 1552
rect 1325 1547 1330 1552
rect 1373 1547 1378 1552
rect 1437 1547 1442 1552
rect 1213 1537 1218 1542
rect 1373 1537 1378 1542
rect 1453 1537 1458 1542
rect 1613 1537 1618 1542
rect 1917 1547 1922 1552
rect 2077 1547 2082 1552
rect 2573 1547 2578 1552
rect 2765 1547 2770 1552
rect 3469 1547 3474 1552
rect 589 1527 594 1532
rect 1229 1527 1234 1532
rect 2477 1537 2482 1542
rect 2253 1527 2258 1532
rect 2789 1527 2794 1532
rect 573 1517 578 1522
rect 1037 1517 1042 1522
rect 2189 1517 2194 1522
rect 365 1507 370 1512
rect 1101 1507 1106 1512
rect 1229 1507 1234 1512
rect 992 1503 994 1507
rect 994 1503 997 1507
rect 1002 1503 1005 1507
rect 1005 1503 1007 1507
rect 992 1502 997 1503
rect 1002 1502 1007 1503
rect 1309 1497 1314 1502
rect 1405 1507 1410 1512
rect 2061 1507 2066 1512
rect 2024 1503 2026 1507
rect 2026 1503 2029 1507
rect 2034 1503 2037 1507
rect 2037 1503 2039 1507
rect 2024 1502 2029 1503
rect 2034 1502 2039 1503
rect 3040 1503 3042 1507
rect 3042 1503 3045 1507
rect 3050 1503 3053 1507
rect 3053 1503 3055 1507
rect 3040 1502 3045 1503
rect 3050 1502 3055 1503
rect 1661 1497 1666 1502
rect 1901 1497 1906 1502
rect 1213 1487 1218 1492
rect 1629 1487 1634 1492
rect 1949 1487 1954 1492
rect 2077 1487 2082 1492
rect 2125 1497 2130 1502
rect 2157 1497 2162 1502
rect 2285 1497 2290 1502
rect 2301 1497 2306 1502
rect 2349 1497 2354 1502
rect 893 1477 898 1482
rect 1325 1477 1330 1482
rect 1917 1477 1922 1482
rect 2493 1487 2498 1492
rect 2653 1487 2658 1492
rect 3325 1477 3330 1482
rect 1021 1467 1026 1472
rect 1261 1467 1266 1472
rect 1277 1467 1282 1472
rect 1213 1457 1218 1462
rect 1629 1467 1634 1472
rect 2013 1467 2018 1472
rect 2045 1467 2050 1472
rect 2349 1467 2354 1472
rect 1389 1457 1394 1462
rect 1421 1457 1426 1462
rect 2317 1457 2322 1462
rect 1117 1447 1122 1452
rect 1837 1447 1842 1452
rect 2429 1447 2434 1452
rect 2461 1447 2466 1452
rect 1469 1437 1474 1442
rect 1613 1437 1618 1442
rect 1709 1437 1714 1442
rect 1757 1437 1762 1442
rect 2381 1437 2386 1442
rect 2573 1437 2578 1442
rect 1485 1427 1490 1432
rect 1565 1427 1570 1432
rect 1885 1427 1890 1432
rect 1933 1427 1938 1432
rect 2077 1427 2082 1432
rect 2397 1427 2402 1432
rect 829 1417 834 1422
rect 845 1417 850 1422
rect 1421 1417 1426 1422
rect 1021 1407 1026 1412
rect 1069 1407 1074 1412
rect 1165 1407 1170 1412
rect 480 1403 482 1407
rect 482 1403 485 1407
rect 490 1403 493 1407
rect 493 1403 495 1407
rect 480 1402 485 1403
rect 490 1402 495 1403
rect 1789 1407 1794 1412
rect 2653 1407 2658 1412
rect 1512 1403 1514 1407
rect 1514 1403 1517 1407
rect 1522 1403 1525 1407
rect 1525 1403 1527 1407
rect 1512 1402 1517 1403
rect 1522 1402 1527 1403
rect 2536 1403 2538 1407
rect 2538 1403 2541 1407
rect 2546 1403 2549 1407
rect 2549 1403 2551 1407
rect 2536 1402 2541 1403
rect 2546 1402 2551 1403
rect 1501 1397 1506 1402
rect 1533 1397 1538 1402
rect 1581 1397 1586 1402
rect 1741 1397 1746 1402
rect 1773 1397 1778 1402
rect 1869 1397 1874 1402
rect 2605 1397 2610 1402
rect 1341 1387 1346 1392
rect 2365 1387 2370 1392
rect 2573 1387 2578 1392
rect 1501 1377 1506 1382
rect 2429 1377 2434 1382
rect 2621 1377 2626 1382
rect 893 1367 898 1372
rect 1325 1367 1330 1372
rect 509 1357 514 1362
rect 1325 1357 1330 1362
rect 1437 1357 1442 1362
rect 1485 1357 1490 1362
rect 1613 1357 1618 1362
rect 1677 1357 1682 1362
rect 1869 1367 1874 1372
rect 2701 1367 2706 1372
rect 2237 1357 2242 1362
rect 2365 1357 2370 1362
rect 973 1347 978 1352
rect 957 1337 962 1342
rect 1389 1347 1394 1352
rect 1101 1337 1106 1342
rect 1149 1337 1154 1342
rect 1325 1337 1330 1342
rect 1581 1347 1586 1352
rect 1597 1347 1602 1352
rect 1693 1347 1698 1352
rect 1709 1347 1714 1352
rect 1949 1347 1954 1352
rect 1997 1347 2002 1352
rect 2173 1347 2178 1352
rect 1597 1337 1602 1342
rect 1661 1337 1666 1342
rect 1885 1337 1890 1342
rect 1981 1337 1986 1342
rect 2093 1337 2098 1342
rect 2237 1337 2242 1342
rect 2365 1337 2370 1342
rect 2525 1337 2530 1342
rect 2573 1337 2578 1342
rect 3485 1337 3490 1342
rect 909 1327 914 1332
rect 1501 1327 1506 1332
rect 2013 1327 2018 1332
rect 2997 1327 3002 1332
rect 973 1317 978 1322
rect 1037 1317 1042 1322
rect 1709 1317 1714 1322
rect 1725 1317 1730 1322
rect 1773 1317 1778 1322
rect 2013 1317 2018 1322
rect 2269 1317 2274 1322
rect 2285 1317 2290 1322
rect 1021 1307 1026 1312
rect 1069 1307 1074 1312
rect 1501 1307 1506 1312
rect 992 1303 994 1307
rect 994 1303 997 1307
rect 1002 1303 1005 1307
rect 1005 1303 1007 1307
rect 992 1302 997 1303
rect 1002 1302 1007 1303
rect 1037 1297 1042 1302
rect 1981 1307 1986 1312
rect 2024 1303 2026 1307
rect 2026 1303 2029 1307
rect 2034 1303 2037 1307
rect 2037 1303 2039 1307
rect 2024 1302 2029 1303
rect 2034 1302 2039 1303
rect 2061 1307 2066 1312
rect 2237 1307 2242 1312
rect 3040 1303 3042 1307
rect 3042 1303 3045 1307
rect 3050 1303 3053 1307
rect 3053 1303 3055 1307
rect 3040 1302 3045 1303
rect 3050 1302 3055 1303
rect 1629 1287 1634 1292
rect 1661 1287 1666 1292
rect 1965 1297 1970 1302
rect 2045 1297 2050 1302
rect 2173 1297 2178 1302
rect 2413 1297 2418 1302
rect 2573 1297 2578 1302
rect 2749 1297 2754 1302
rect 2077 1287 2082 1292
rect 2093 1287 2098 1292
rect 2205 1287 2210 1292
rect 957 1277 962 1282
rect 1133 1277 1138 1282
rect 781 1267 786 1272
rect 1021 1267 1026 1272
rect 1293 1267 1298 1272
rect 1405 1277 1410 1282
rect 1053 1257 1058 1262
rect 1309 1257 1314 1262
rect 1325 1257 1330 1262
rect 1421 1267 1426 1272
rect 1677 1267 1682 1272
rect 2301 1277 2306 1282
rect 2413 1267 2418 1272
rect 2445 1267 2450 1272
rect 2509 1267 2514 1272
rect 2637 1267 2642 1272
rect 1357 1257 1362 1262
rect 1437 1257 1442 1262
rect 1085 1247 1090 1252
rect 2589 1257 2594 1262
rect 2157 1247 2162 1252
rect 2237 1247 2242 1252
rect 1197 1237 1202 1242
rect 2317 1237 2322 1242
rect 2829 1237 2834 1242
rect 1597 1227 1602 1232
rect 1693 1227 1698 1232
rect 1741 1227 1746 1232
rect 2573 1227 2578 1232
rect 2077 1217 2082 1222
rect 949 1207 954 1212
rect 973 1207 978 1212
rect 1645 1207 1650 1212
rect 2621 1207 2626 1212
rect 2685 1207 2690 1212
rect 480 1203 482 1207
rect 482 1203 485 1207
rect 490 1203 493 1207
rect 493 1203 495 1207
rect 480 1202 485 1203
rect 490 1202 495 1203
rect 1512 1203 1514 1207
rect 1514 1203 1517 1207
rect 1522 1203 1525 1207
rect 1525 1203 1527 1207
rect 1512 1202 1517 1203
rect 1522 1202 1527 1203
rect 2536 1203 2538 1207
rect 2538 1203 2541 1207
rect 2546 1203 2549 1207
rect 2549 1203 2551 1207
rect 2536 1202 2541 1203
rect 2546 1202 2551 1203
rect 941 1197 946 1202
rect 1533 1197 1538 1202
rect 2077 1197 2082 1202
rect 1325 1187 1330 1192
rect 1389 1187 1394 1192
rect 1101 1177 1106 1182
rect 1229 1177 1234 1182
rect 1245 1177 1250 1182
rect 2093 1177 2098 1182
rect 461 1167 466 1172
rect 1325 1167 1330 1172
rect 1341 1167 1346 1172
rect 1485 1167 1490 1172
rect 1581 1167 1586 1172
rect 1277 1157 1282 1162
rect 1325 1157 1330 1162
rect 1709 1157 1714 1162
rect 1757 1157 1762 1162
rect 2429 1167 2434 1172
rect 749 1147 754 1152
rect 1037 1147 1042 1152
rect 1133 1147 1138 1152
rect 1373 1147 1378 1152
rect 1581 1147 1586 1152
rect 1869 1147 1874 1152
rect 1965 1147 1970 1152
rect 2109 1147 2114 1152
rect 2237 1147 2242 1152
rect 1181 1137 1186 1142
rect 1277 1137 1282 1142
rect 1309 1137 1314 1142
rect 1373 1137 1378 1142
rect 1645 1137 1650 1142
rect 2605 1137 2610 1142
rect 669 1127 674 1132
rect 861 1127 866 1132
rect 1181 1117 1186 1122
rect 1565 1127 1570 1132
rect 1597 1127 1602 1132
rect 2061 1127 2066 1132
rect 2557 1127 2562 1132
rect 1421 1118 1422 1122
rect 1422 1118 1426 1122
rect 1421 1117 1426 1118
rect 1645 1117 1650 1122
rect 1677 1117 1682 1122
rect 1709 1117 1714 1122
rect 1261 1107 1266 1112
rect 1325 1107 1330 1112
rect 1341 1107 1346 1112
rect 1453 1107 1458 1112
rect 1645 1107 1650 1112
rect 1677 1107 1682 1112
rect 992 1103 994 1107
rect 994 1103 997 1107
rect 1002 1103 1005 1107
rect 1005 1103 1007 1107
rect 992 1102 997 1103
rect 1002 1102 1007 1103
rect 925 1097 930 1102
rect 1037 1097 1042 1102
rect 1197 1097 1202 1102
rect 1709 1097 1714 1102
rect 1949 1107 1954 1112
rect 2077 1107 2082 1112
rect 2024 1103 2026 1107
rect 2026 1103 2029 1107
rect 2034 1103 2037 1107
rect 2037 1103 2039 1107
rect 2024 1102 2029 1103
rect 2034 1102 2039 1103
rect 3040 1103 3042 1107
rect 3042 1103 3045 1107
rect 3050 1103 3053 1107
rect 3053 1103 3055 1107
rect 3040 1102 3045 1103
rect 3050 1102 3055 1103
rect 2045 1097 2050 1102
rect 2413 1097 2418 1102
rect 1149 1087 1154 1092
rect 1341 1087 1346 1092
rect 1405 1087 1410 1092
rect 1437 1087 1442 1092
rect 1773 1087 1778 1092
rect 2285 1087 2290 1092
rect 2653 1087 2658 1092
rect 1165 1077 1170 1082
rect 1597 1077 1602 1082
rect 1837 1077 1842 1082
rect 2397 1077 2402 1082
rect 957 1067 962 1072
rect 1469 1067 1474 1072
rect 1485 1067 1490 1072
rect 1741 1067 1746 1072
rect 1805 1067 1810 1072
rect 2013 1067 2018 1072
rect 2861 1067 2866 1072
rect 1117 1057 1122 1062
rect 1853 1057 1858 1062
rect 2349 1057 2354 1062
rect 877 1047 882 1052
rect 973 1047 978 1052
rect 1213 1047 1218 1052
rect 1613 1037 1618 1042
rect 1741 1037 1746 1042
rect 1981 1037 1986 1042
rect 733 1027 738 1032
rect 877 1027 882 1032
rect 2109 1027 2114 1032
rect 2205 1027 2210 1032
rect 797 1017 802 1022
rect 1245 1017 1250 1022
rect 1277 1017 1282 1022
rect 1341 1017 1346 1022
rect 941 1007 946 1012
rect 1493 1007 1498 1012
rect 480 1003 482 1007
rect 482 1003 485 1007
rect 490 1003 493 1007
rect 493 1003 495 1007
rect 480 1002 485 1003
rect 490 1002 495 1003
rect 1512 1003 1514 1007
rect 1514 1003 1517 1007
rect 1522 1003 1525 1007
rect 1525 1003 1527 1007
rect 1512 1002 1517 1003
rect 1522 1002 1527 1003
rect 1741 1007 1746 1012
rect 2536 1003 2538 1007
rect 2538 1003 2541 1007
rect 2546 1003 2549 1007
rect 2549 1003 2551 1007
rect 2536 1002 2541 1003
rect 2546 1002 2551 1003
rect 829 997 834 1002
rect 1069 998 1070 1002
rect 1070 998 1074 1002
rect 1069 997 1074 998
rect 1581 997 1586 1002
rect 1981 997 1986 1002
rect 1213 987 1218 992
rect 1229 987 1234 992
rect 1245 977 1250 982
rect 1261 987 1266 992
rect 1277 987 1282 992
rect 1693 987 1698 992
rect 3517 987 3522 992
rect 1469 977 1474 982
rect 1933 977 1938 982
rect 1949 977 1954 982
rect 2013 977 2018 982
rect 1469 957 1474 962
rect 1645 957 1650 962
rect 2045 957 2050 962
rect 2125 957 2130 962
rect 2205 957 2210 962
rect 957 937 962 942
rect 1757 947 1762 952
rect 1293 937 1298 942
rect 1469 937 1474 942
rect 1485 937 1490 942
rect 1933 937 1938 942
rect 2685 937 2690 942
rect 1325 927 1330 932
rect 1789 927 1794 932
rect 2445 927 2450 932
rect 701 917 706 922
rect 1357 917 1362 922
rect 1709 917 1714 922
rect 1021 907 1026 912
rect 1293 907 1298 912
rect 1677 907 1682 912
rect 2013 907 2018 912
rect 2077 907 2082 912
rect 2093 907 2098 912
rect 992 903 994 907
rect 994 903 997 907
rect 1002 903 1005 907
rect 1005 903 1007 907
rect 992 902 997 903
rect 1002 902 1007 903
rect 2024 903 2026 907
rect 2026 903 2029 907
rect 2034 903 2037 907
rect 2037 903 2039 907
rect 2024 902 2029 903
rect 2034 902 2039 903
rect 3040 903 3042 907
rect 3042 903 3045 907
rect 3050 903 3053 907
rect 3053 903 3055 907
rect 3040 902 3045 903
rect 3050 902 3055 903
rect 1213 897 1218 902
rect 1405 897 1410 902
rect 1245 887 1250 892
rect 1565 887 1570 892
rect 1581 887 1586 892
rect 1725 887 1730 892
rect 1917 897 1922 902
rect 2045 897 2050 902
rect 2845 887 2850 892
rect 1181 877 1186 882
rect 813 867 818 872
rect 1245 867 1250 872
rect 1485 867 1490 872
rect 877 857 882 862
rect 1053 857 1058 862
rect 1485 857 1490 862
rect 1429 847 1434 852
rect 1645 847 1650 852
rect 717 837 722 842
rect 1309 827 1314 832
rect 480 803 482 807
rect 482 803 485 807
rect 490 803 493 807
rect 493 803 495 807
rect 480 802 485 803
rect 490 802 495 803
rect 797 797 802 802
rect 1565 807 1570 812
rect 1512 803 1514 807
rect 1514 803 1517 807
rect 1522 803 1525 807
rect 1525 803 1527 807
rect 1512 802 1517 803
rect 1522 802 1527 803
rect 2536 803 2538 807
rect 2538 803 2541 807
rect 2546 803 2549 807
rect 2549 803 2551 807
rect 2536 802 2541 803
rect 2546 802 2551 803
rect 1181 797 1186 802
rect 2093 797 2098 802
rect 1165 787 1170 792
rect 1253 767 1258 772
rect 973 757 978 762
rect 1181 757 1186 762
rect 1309 757 1314 762
rect 2701 767 2706 772
rect 1389 757 1394 762
rect 1997 757 2002 762
rect 2749 757 2754 762
rect 781 747 786 752
rect 1725 747 1730 752
rect 1117 737 1122 742
rect 1741 747 1746 752
rect 909 727 914 732
rect 925 727 930 732
rect 1277 727 1282 732
rect 1997 727 2002 732
rect 2301 727 2306 732
rect 669 717 674 722
rect 1485 707 1490 712
rect 992 703 994 707
rect 994 703 997 707
rect 1002 703 1005 707
rect 1005 703 1007 707
rect 992 702 997 703
rect 1002 702 1007 703
rect 2024 703 2026 707
rect 2026 703 2029 707
rect 2034 703 2037 707
rect 2037 703 2039 707
rect 2024 702 2029 703
rect 2034 702 2039 703
rect 3040 703 3042 707
rect 3042 703 3045 707
rect 3050 703 3053 707
rect 3053 703 3055 707
rect 3040 702 3045 703
rect 3050 702 3055 703
rect 365 697 370 702
rect 893 697 898 702
rect 1405 697 1410 702
rect 1533 697 1538 702
rect 1693 697 1698 702
rect 1501 687 1506 692
rect 1709 687 1714 692
rect 1085 677 1090 682
rect 1245 677 1250 682
rect 1277 677 1282 682
rect 1501 677 1506 682
rect 2045 677 2050 682
rect 2173 677 2178 682
rect 509 667 514 672
rect 1341 667 1346 672
rect 717 657 722 662
rect 1277 657 1282 662
rect 1693 657 1698 662
rect 1933 657 1938 662
rect 605 637 610 642
rect 1245 647 1250 652
rect 1485 647 1490 652
rect 1501 647 1506 652
rect 1325 637 1330 642
rect 749 627 754 632
rect 1101 627 1106 632
rect 1309 627 1314 632
rect 685 617 690 622
rect 877 617 882 622
rect 1549 617 1554 622
rect 861 607 866 612
rect 1037 607 1042 612
rect 480 603 482 607
rect 482 603 485 607
rect 490 603 493 607
rect 493 603 495 607
rect 480 602 485 603
rect 490 602 495 603
rect 1512 603 1514 607
rect 1514 603 1517 607
rect 1522 603 1525 607
rect 1525 603 1527 607
rect 1512 602 1517 603
rect 1522 602 1527 603
rect 2536 603 2538 607
rect 2538 603 2541 607
rect 2546 603 2549 607
rect 2549 603 2551 607
rect 2536 602 2541 603
rect 2546 602 2551 603
rect 797 587 802 592
rect 877 587 882 592
rect 893 587 898 592
rect 1101 587 1106 592
rect 1405 577 1410 582
rect 1661 577 1666 582
rect 1133 557 1138 562
rect 1821 557 1826 562
rect 925 547 930 552
rect 973 547 978 552
rect 1117 547 1122 552
rect 1405 547 1410 552
rect 2221 537 2226 542
rect 1373 517 1378 522
rect 2141 517 2146 522
rect 1949 507 1954 512
rect 992 503 994 507
rect 994 503 997 507
rect 1002 503 1005 507
rect 1005 503 1007 507
rect 992 502 997 503
rect 1002 502 1007 503
rect 2024 503 2026 507
rect 2026 503 2029 507
rect 2034 503 2037 507
rect 2037 503 2039 507
rect 2024 502 2029 503
rect 2034 502 2039 503
rect 3040 503 3042 507
rect 3042 503 3045 507
rect 3050 503 3053 507
rect 3053 503 3055 507
rect 3040 502 3045 503
rect 3050 502 3055 503
rect 973 497 978 502
rect 1021 497 1026 502
rect 2221 477 2226 482
rect 1341 467 1346 472
rect 813 457 818 462
rect 2685 457 2690 462
rect 1133 437 1138 442
rect 1021 417 1026 422
rect 1037 417 1042 422
rect 2077 417 2082 422
rect 480 403 482 407
rect 482 403 485 407
rect 490 403 493 407
rect 493 403 495 407
rect 480 402 485 403
rect 490 402 495 403
rect 1512 403 1514 407
rect 1514 403 1517 407
rect 1522 403 1525 407
rect 1525 403 1527 407
rect 1512 402 1517 403
rect 1522 402 1527 403
rect 2536 403 2538 407
rect 2538 403 2541 407
rect 2546 403 2549 407
rect 2549 403 2551 407
rect 2536 402 2541 403
rect 2546 402 2551 403
rect 3437 377 3442 382
rect 589 347 594 352
rect 541 337 546 342
rect 621 328 622 332
rect 622 328 626 332
rect 621 327 626 328
rect 637 327 642 332
rect 669 327 674 332
rect 2765 317 2770 322
rect 992 303 994 307
rect 994 303 997 307
rect 1002 303 1005 307
rect 1005 303 1007 307
rect 992 302 997 303
rect 1002 302 1007 303
rect 2024 303 2026 307
rect 2026 303 2029 307
rect 2034 303 2037 307
rect 2037 303 2039 307
rect 2024 302 2029 303
rect 2034 302 2039 303
rect 3040 303 3042 307
rect 3042 303 3045 307
rect 3050 303 3053 307
rect 3053 303 3055 307
rect 3040 302 3045 303
rect 3050 302 3055 303
rect 2621 257 2626 262
rect 480 203 482 207
rect 482 203 485 207
rect 490 203 493 207
rect 493 203 495 207
rect 480 202 485 203
rect 490 202 495 203
rect 1512 203 1514 207
rect 1514 203 1517 207
rect 1522 203 1525 207
rect 1525 203 1527 207
rect 1512 202 1517 203
rect 1522 202 1527 203
rect 2536 203 2538 207
rect 2538 203 2541 207
rect 2546 203 2549 207
rect 2549 203 2551 207
rect 2536 202 2541 203
rect 2546 202 2551 203
rect 701 187 706 192
rect 992 103 994 107
rect 994 103 997 107
rect 1002 103 1005 107
rect 1005 103 1007 107
rect 992 102 997 103
rect 1002 102 1007 103
rect 2024 103 2026 107
rect 2026 103 2029 107
rect 2034 103 2037 107
rect 2037 103 2039 107
rect 2024 102 2029 103
rect 2034 102 2039 103
rect 3040 103 3042 107
rect 3042 103 3045 107
rect 3050 103 3053 107
rect 3053 103 3055 107
rect 3040 102 3045 103
rect 3050 102 3055 103
rect 605 77 610 82
rect 3485 77 3490 82
rect 3325 67 3330 72
rect 3357 67 3362 72
rect 2765 17 2770 22
rect 480 3 482 7
rect 482 3 485 7
rect 490 3 493 7
rect 493 3 495 7
rect 480 2 485 3
rect 490 2 495 3
rect 1512 3 1514 7
rect 1514 3 1517 7
rect 1522 3 1525 7
rect 1525 3 1527 7
rect 1512 2 1517 3
rect 1522 2 1527 3
rect 2536 3 2538 7
rect 2538 3 2541 7
rect 2546 3 2549 7
rect 2549 3 2551 7
rect 2536 2 2541 3
rect 2546 2 2551 3
<< metal6 >>
rect 480 3207 496 3330
rect 485 3202 490 3207
rect 495 3202 496 3207
rect 480 3007 496 3202
rect 485 3002 490 3007
rect 495 3002 496 3007
rect 480 2807 496 3002
rect 485 2802 490 2807
rect 495 2802 496 2807
rect 480 2607 496 2802
rect 485 2602 490 2607
rect 495 2602 496 2607
rect 480 2407 496 2602
rect 485 2402 490 2407
rect 495 2402 496 2407
rect 480 2207 496 2402
rect 992 3307 1008 3330
rect 997 3302 1002 3307
rect 1007 3302 1008 3307
rect 992 3107 1008 3302
rect 997 3102 1002 3107
rect 1007 3102 1008 3107
rect 992 2907 1008 3102
rect 997 2902 1002 2907
rect 1007 2902 1008 2907
rect 992 2707 1008 2902
rect 997 2702 1002 2707
rect 1007 2702 1008 2707
rect 992 2507 1008 2702
rect 1053 2542 1058 3227
rect 1133 2552 1138 3297
rect 1512 3207 1528 3330
rect 1517 3202 1522 3207
rect 1527 3202 1528 3207
rect 1512 3007 1528 3202
rect 2024 3307 2040 3330
rect 2029 3302 2034 3307
rect 2039 3302 2040 3307
rect 2024 3107 2040 3302
rect 2029 3102 2034 3107
rect 2039 3102 2040 3107
rect 1517 3002 1522 3007
rect 1527 3002 1528 3007
rect 1512 2807 1528 3002
rect 1517 2802 1522 2807
rect 1527 2802 1528 2807
rect 1512 2607 1528 2802
rect 1517 2602 1522 2607
rect 1527 2602 1528 2607
rect 997 2502 1002 2507
rect 1007 2502 1008 2507
rect 485 2202 490 2207
rect 495 2202 496 2207
rect 480 2007 496 2202
rect 485 2002 490 2007
rect 495 2002 496 2007
rect 480 1807 496 2002
rect 485 1802 490 1807
rect 495 1802 496 1807
rect 365 702 370 1507
rect 461 1172 466 1727
rect 480 1607 496 1802
rect 485 1602 490 1607
rect 495 1602 496 1607
rect 480 1407 496 1602
rect 485 1402 490 1407
rect 495 1402 496 1407
rect 480 1207 496 1402
rect 541 2222 546 2337
rect 485 1202 490 1207
rect 495 1202 496 1207
rect 480 1007 496 1202
rect 485 1002 490 1007
rect 495 1002 496 1007
rect 480 807 496 1002
rect 485 802 490 807
rect 495 802 496 807
rect 480 607 496 802
rect 509 672 514 1357
rect 485 602 490 607
rect 495 602 496 607
rect 480 407 496 602
rect 485 402 490 407
rect 495 402 496 407
rect 480 207 496 402
rect 541 342 546 2217
rect 557 1702 562 2257
rect 573 1522 578 1867
rect 589 1532 594 2017
rect 605 1602 610 2167
rect 717 2132 722 2307
rect 621 1682 626 1837
rect 589 352 594 1527
rect 485 202 490 207
rect 495 202 496 207
rect 480 7 496 202
rect 605 82 610 637
rect 621 332 626 1657
rect 637 332 642 1867
rect 669 1132 674 1697
rect 669 722 674 1127
rect 669 332 674 717
rect 685 622 690 1827
rect 717 1542 722 2127
rect 992 2307 1008 2502
rect 997 2302 1002 2307
rect 1007 2302 1008 2307
rect 992 2107 1008 2302
rect 1512 2407 1528 2602
rect 1533 2412 1538 2517
rect 1517 2402 1522 2407
rect 1527 2402 1528 2407
rect 1501 2192 1506 2207
rect 1512 2207 1528 2402
rect 1517 2202 1522 2207
rect 1527 2202 1528 2207
rect 997 2102 1002 2107
rect 1007 2102 1008 2107
rect 845 2007 853 2012
rect 733 1032 738 1997
rect 749 1802 754 1827
rect 701 192 706 917
rect 717 662 722 837
rect 749 632 754 1147
rect 781 752 786 1267
rect 797 1022 802 1627
rect 845 1422 850 2007
rect 829 1002 834 1417
rect 797 592 802 797
rect 813 462 818 867
rect 861 612 866 1127
rect 877 1052 882 1597
rect 893 1482 898 1917
rect 992 1907 1008 2102
rect 997 1902 1002 1907
rect 1007 1902 1008 1907
rect 909 1812 914 1897
rect 877 862 882 1027
rect 893 702 898 1367
rect 909 1332 914 1807
rect 957 1772 962 1797
rect 909 732 914 1327
rect 925 1102 930 1727
rect 941 1212 946 1657
rect 957 1652 962 1717
rect 973 1352 978 1867
rect 992 1707 1008 1902
rect 997 1702 1002 1707
rect 1007 1702 1008 1707
rect 992 1507 1008 1702
rect 997 1502 1002 1507
rect 1007 1502 1008 1507
rect 957 1282 962 1337
rect 973 1212 978 1317
rect 941 1207 949 1212
rect 992 1307 1008 1502
rect 1021 1472 1026 1697
rect 1037 1522 1042 1977
rect 1021 1457 1026 1467
rect 1021 1312 1026 1407
rect 997 1302 1002 1307
rect 1007 1302 1008 1307
rect 941 1012 946 1197
rect 992 1107 1008 1302
rect 1037 1302 1042 1317
rect 997 1102 1002 1107
rect 1007 1102 1008 1107
rect 957 942 962 1067
rect 973 762 978 1047
rect 992 907 1008 1102
rect 1021 912 1026 1267
rect 1053 1262 1058 1857
rect 1069 1412 1074 1807
rect 1085 1602 1090 1727
rect 1101 1512 1106 1897
rect 1165 1842 1170 1857
rect 1341 1827 1349 1832
rect 1181 1652 1186 1657
rect 1130 1647 1186 1652
rect 1117 1552 1122 1617
rect 1229 1592 1234 1787
rect 1149 1562 1154 1577
rect 1037 1102 1042 1147
rect 997 902 1002 907
rect 1007 902 1008 907
rect 877 592 882 617
rect 893 592 898 697
rect 925 552 930 727
rect 992 707 1008 902
rect 1053 862 1058 1257
rect 1069 1002 1074 1307
rect 997 702 1002 707
rect 1007 702 1008 707
rect 973 502 978 547
rect 992 507 1008 702
rect 1085 682 1090 1247
rect 1101 1182 1106 1337
rect 1117 1062 1122 1447
rect 1165 1412 1170 1587
rect 1133 1152 1138 1277
rect 1149 1092 1154 1337
rect 1181 1142 1186 1547
rect 1213 1492 1218 1537
rect 1229 1512 1234 1527
rect 1261 1472 1266 1737
rect 1309 1662 1314 1707
rect 1277 1652 1282 1657
rect 1277 1647 1301 1652
rect 1165 792 1170 1077
rect 1181 882 1186 1117
rect 1197 1102 1202 1237
rect 1213 1052 1218 1457
rect 1229 992 1234 1177
rect 1245 1022 1250 1177
rect 1277 1162 1282 1467
rect 1293 1272 1298 1567
rect 1309 1552 1314 1587
rect 1325 1552 1330 1747
rect 1309 1262 1314 1497
rect 1325 1372 1330 1477
rect 1341 1392 1346 1827
rect 1373 1552 1378 1767
rect 1405 1732 1410 2057
rect 1512 2007 1528 2202
rect 1709 2192 1714 2327
rect 1725 2272 1730 3057
rect 1789 2927 1797 2932
rect 1517 2002 1522 2007
rect 1527 2002 1528 2007
rect 1421 1732 1426 1777
rect 1389 1612 1394 1657
rect 1389 1607 1426 1612
rect 1421 1582 1426 1607
rect 1325 1342 1330 1357
rect 1325 1262 1330 1337
rect 1325 1172 1330 1187
rect 1261 992 1266 1107
rect 1277 1022 1282 1137
rect 1213 902 1218 987
rect 1245 892 1250 977
rect 1181 762 1186 797
rect 1245 772 1250 867
rect 1245 767 1253 772
rect 997 502 1002 507
rect 1007 502 1008 507
rect 992 307 1008 502
rect 1021 422 1026 497
rect 1037 422 1042 607
rect 1101 592 1106 627
rect 1117 552 1122 737
rect 1277 732 1282 987
rect 1293 912 1298 937
rect 1309 832 1314 1137
rect 1325 1112 1330 1157
rect 1341 1112 1346 1167
rect 1341 1022 1346 1087
rect 1245 652 1250 677
rect 1277 662 1282 677
rect 1309 632 1314 757
rect 1325 642 1330 927
rect 1357 922 1362 1257
rect 1373 1152 1378 1537
rect 1389 1462 1394 1567
rect 1405 1512 1410 1577
rect 1437 1572 1442 1747
rect 1389 1352 1394 1457
rect 1421 1422 1426 1457
rect 1437 1362 1442 1547
rect 1133 442 1138 557
rect 1341 472 1346 667
rect 1373 522 1378 1137
rect 1389 762 1394 1187
rect 1405 1092 1410 1277
rect 1421 1122 1426 1267
rect 1437 1092 1442 1257
rect 1453 1112 1458 1537
rect 1469 1442 1474 1827
rect 1485 1782 1490 1837
rect 1501 1602 1506 1847
rect 1512 1807 1528 2002
rect 1517 1802 1522 1807
rect 1527 1802 1528 1807
rect 1512 1607 1528 1802
rect 1517 1602 1522 1607
rect 1527 1602 1528 1607
rect 1485 1362 1490 1427
rect 1512 1407 1528 1602
rect 1517 1402 1522 1407
rect 1527 1402 1528 1407
rect 1501 1382 1506 1397
rect 1501 1312 1506 1327
rect 1512 1207 1528 1402
rect 1533 1402 1538 2167
rect 1789 2132 1794 2927
rect 1821 2922 1826 2937
rect 2024 2907 2040 3102
rect 2536 3207 2552 3330
rect 2541 3202 2546 3207
rect 2551 3202 2552 3207
rect 2029 2902 2034 2907
rect 2039 2902 2040 2907
rect 1997 2612 2002 2867
rect 2024 2707 2040 2902
rect 2029 2702 2034 2707
rect 2039 2702 2040 2707
rect 2024 2507 2040 2702
rect 2029 2502 2034 2507
rect 2039 2502 2040 2507
rect 2024 2307 2040 2502
rect 2029 2302 2034 2307
rect 2039 2302 2040 2307
rect 2024 2107 2040 2302
rect 2029 2102 2034 2107
rect 2039 2102 2040 2107
rect 1581 1672 1586 2067
rect 1549 1607 1557 1612
rect 1517 1202 1522 1207
rect 1527 1202 1528 1207
rect 1485 1072 1490 1167
rect 1469 982 1474 1067
rect 1498 1007 1506 1012
rect 1469 942 1474 957
rect 1405 702 1410 897
rect 1485 872 1490 937
rect 1485 852 1490 857
rect 1434 847 1490 852
rect 1485 652 1490 707
rect 1501 692 1506 1007
rect 1512 1007 1528 1202
rect 1517 1002 1522 1007
rect 1527 1002 1528 1007
rect 1512 807 1528 1002
rect 1517 802 1522 807
rect 1527 802 1528 807
rect 1501 652 1506 677
rect 1512 607 1528 802
rect 1533 702 1538 1197
rect 1549 622 1554 1607
rect 1565 1132 1570 1427
rect 1581 1352 1586 1397
rect 1597 1352 1602 1917
rect 1613 1442 1618 1537
rect 1629 1492 1634 1967
rect 1597 1232 1602 1337
rect 1581 1152 1586 1167
rect 1597 1082 1602 1127
rect 1613 1042 1618 1357
rect 1629 1292 1634 1467
rect 1645 1212 1650 2007
rect 1661 1692 1666 1967
rect 1677 1872 1682 2017
rect 1661 1342 1666 1497
rect 1677 1362 1682 1767
rect 1693 1352 1698 1877
rect 1709 1782 1714 1877
rect 1725 1782 1730 1857
rect 1709 1582 1714 1687
rect 1725 1612 1730 1767
rect 1709 1352 1714 1437
rect 1741 1402 1746 2057
rect 1773 1922 1778 2017
rect 1757 1842 1762 1897
rect 1757 1602 1762 1667
rect 1757 1442 1762 1587
rect 1773 1402 1778 1897
rect 1789 1672 1794 1927
rect 1645 1122 1650 1137
rect 1581 892 1586 997
rect 1645 962 1650 1107
rect 1565 812 1570 887
rect 1645 852 1650 957
rect 1517 602 1522 607
rect 1527 602 1528 607
rect 1405 552 1410 577
rect 997 302 1002 307
rect 1007 302 1008 307
rect 992 107 1008 302
rect 997 102 1002 107
rect 1007 102 1008 107
rect 485 2 490 7
rect 495 2 496 7
rect 480 -30 496 2
rect 992 -30 1008 102
rect 1512 407 1528 602
rect 1661 582 1666 1287
rect 1677 1122 1682 1267
rect 1677 912 1682 1107
rect 1693 992 1698 1227
rect 1709 1162 1714 1317
rect 1709 1102 1714 1117
rect 1693 662 1698 697
rect 1709 692 1714 917
rect 1725 892 1730 1317
rect 1741 1072 1746 1227
rect 1741 1012 1746 1037
rect 1757 952 1762 1157
rect 1773 1092 1778 1317
rect 1789 932 1794 1407
rect 1805 1072 1810 1687
rect 1730 747 1741 752
rect 1821 562 1826 1717
rect 1837 1672 1842 2047
rect 1853 1592 1858 1667
rect 1885 1592 1890 1837
rect 1837 1082 1842 1447
rect 1853 1062 1858 1557
rect 1869 1402 1874 1587
rect 1901 1502 1906 1967
rect 1949 1952 1954 1977
rect 1917 1552 1922 1947
rect 1933 1582 1938 1917
rect 1997 1832 2002 2007
rect 2024 1907 2040 2102
rect 2029 1902 2034 1907
rect 2039 1902 2040 1907
rect 1949 1492 1954 1717
rect 1869 1152 1874 1367
rect 1885 1342 1890 1427
rect 1917 902 1922 1477
rect 1933 982 1938 1427
rect 1949 1112 1954 1347
rect 1981 1342 1986 1587
rect 1997 1352 2002 1657
rect 2013 1562 2018 1837
rect 2024 1707 2040 1902
rect 2029 1702 2034 1707
rect 2039 1702 2040 1707
rect 2024 1507 2040 1702
rect 2029 1502 2034 1507
rect 2039 1502 2040 1507
rect 2013 1332 2018 1467
rect 1965 1152 1970 1297
rect 1981 1042 1986 1307
rect 2013 1072 2018 1317
rect 2024 1307 2040 1502
rect 2045 1472 2050 2727
rect 2061 1832 2066 2227
rect 2205 2102 2210 2547
rect 2061 1672 2066 1807
rect 2061 1512 2066 1567
rect 2077 1552 2082 1947
rect 2077 1432 2082 1487
rect 2093 1342 2098 1947
rect 2109 1722 2114 1787
rect 2125 1502 2130 1907
rect 2157 1832 2162 1877
rect 2029 1302 2034 1307
rect 2039 1302 2040 1307
rect 2024 1107 2040 1302
rect 2029 1102 2034 1107
rect 2039 1102 2040 1107
rect 1981 1002 1986 1037
rect 1933 662 1938 937
rect 1949 512 1954 977
rect 2013 912 2018 977
rect 2024 907 2040 1102
rect 2045 1102 2050 1297
rect 2061 1132 2066 1307
rect 2077 1222 2082 1287
rect 2077 1112 2082 1197
rect 2093 1182 2098 1287
rect 2045 962 2050 1097
rect 2109 1032 2114 1147
rect 2125 962 2130 1497
rect 2029 902 2034 907
rect 2039 902 2040 907
rect 1997 732 2002 757
rect 2024 707 2040 902
rect 2029 702 2034 707
rect 2039 702 2040 707
rect 2024 507 2040 702
rect 2045 682 2050 897
rect 1517 402 1522 407
rect 1527 402 1528 407
rect 1512 207 1528 402
rect 1517 202 1522 207
rect 1527 202 1528 207
rect 1512 7 1528 202
rect 1517 2 1522 7
rect 1527 2 1528 7
rect 1512 -30 1528 2
rect 2029 502 2034 507
rect 2039 502 2040 507
rect 2024 307 2040 502
rect 2077 422 2082 907
rect 2093 802 2098 907
rect 2141 522 2146 1597
rect 2157 1252 2162 1497
rect 2173 1352 2178 2057
rect 2301 1947 2309 1952
rect 2189 1522 2194 1867
rect 2173 682 2178 1297
rect 2205 1292 2210 1687
rect 2205 962 2210 1027
rect 2221 542 2226 1927
rect 2237 1362 2242 1907
rect 2253 1532 2258 1887
rect 2237 1312 2242 1337
rect 2269 1322 2274 1817
rect 2285 1742 2290 1867
rect 2285 1502 2290 1737
rect 2301 1502 2306 1947
rect 2349 1832 2354 1887
rect 2365 1682 2370 1727
rect 2349 1502 2354 1677
rect 2237 1152 2242 1247
rect 2285 1092 2290 1317
rect 2301 732 2306 1277
rect 2317 1242 2322 1457
rect 2349 1062 2354 1467
rect 2365 1392 2370 1607
rect 2381 1442 2386 2107
rect 2397 1712 2402 3087
rect 2536 3007 2552 3202
rect 2541 3002 2546 3007
rect 2551 3002 2552 3007
rect 2365 1342 2370 1357
rect 2397 1082 2402 1427
rect 2413 1302 2418 1797
rect 2429 1452 2434 2077
rect 2461 1452 2466 2507
rect 2477 1742 2482 1837
rect 2477 1542 2482 1567
rect 2493 1492 2498 2327
rect 2413 1102 2418 1267
rect 2429 1172 2434 1377
rect 2509 1272 2514 2207
rect 2525 1792 2530 2877
rect 2536 2807 2552 3002
rect 2541 2802 2546 2807
rect 2551 2802 2552 2807
rect 2536 2607 2552 2802
rect 3040 3307 3056 3330
rect 3045 3302 3050 3307
rect 3055 3302 3056 3307
rect 3040 3107 3056 3302
rect 3045 3102 3050 3107
rect 3055 3102 3056 3107
rect 3040 2907 3056 3102
rect 3045 2902 3050 2907
rect 3055 2902 3056 2907
rect 2541 2602 2546 2607
rect 2551 2602 2552 2607
rect 2536 2407 2552 2602
rect 2541 2402 2546 2407
rect 2551 2402 2552 2407
rect 2536 2207 2552 2402
rect 2541 2202 2546 2207
rect 2551 2202 2552 2207
rect 2536 2007 2552 2202
rect 2541 2002 2546 2007
rect 2551 2002 2552 2007
rect 2536 1807 2552 2002
rect 2541 1802 2546 1807
rect 2551 1802 2552 1807
rect 2525 1342 2530 1747
rect 2536 1607 2552 1802
rect 2541 1602 2546 1607
rect 2551 1602 2552 1607
rect 2536 1407 2552 1602
rect 2541 1402 2546 1407
rect 2551 1402 2552 1407
rect 2445 932 2450 1267
rect 2536 1207 2552 1402
rect 2541 1202 2546 1207
rect 2551 1202 2552 1207
rect 2536 1007 2552 1202
rect 2557 1132 2562 1597
rect 2573 1442 2578 1547
rect 2573 1342 2578 1387
rect 2573 1232 2578 1297
rect 2589 1262 2594 2547
rect 2605 1142 2610 1397
rect 2621 1382 2626 1717
rect 2637 1272 2642 1877
rect 2653 1492 2658 1917
rect 2541 1002 2546 1007
rect 2551 1002 2552 1007
rect 2536 807 2552 1002
rect 2541 802 2546 807
rect 2551 802 2552 807
rect 2221 482 2226 537
rect 2536 607 2552 802
rect 2541 602 2546 607
rect 2551 602 2552 607
rect 2029 302 2034 307
rect 2039 302 2040 307
rect 2024 107 2040 302
rect 2029 102 2034 107
rect 2039 102 2040 107
rect 2024 -30 2040 102
rect 2536 407 2552 602
rect 2541 402 2546 407
rect 2551 402 2552 407
rect 2536 207 2552 402
rect 2621 262 2626 1207
rect 2653 1092 2658 1407
rect 2685 1212 2690 1877
rect 2765 1552 2770 2657
rect 2797 1532 2802 1957
rect 2794 1527 2802 1532
rect 2685 462 2690 937
rect 2701 772 2706 1367
rect 2749 762 2754 1297
rect 2829 1242 2834 1877
rect 2845 892 2850 1847
rect 2861 1072 2866 2737
rect 3040 2707 3056 2902
rect 3045 2702 3050 2707
rect 3055 2702 3056 2707
rect 3040 2507 3056 2702
rect 3045 2502 3050 2507
rect 3055 2502 3056 2507
rect 3040 2307 3056 2502
rect 3045 2302 3050 2307
rect 3055 2302 3056 2307
rect 3040 2107 3056 2302
rect 3373 2302 3378 3007
rect 3045 2102 3050 2107
rect 3055 2102 3056 2107
rect 3040 1907 3056 2102
rect 3045 1902 3050 1907
rect 3055 1902 3056 1907
rect 3005 1332 3010 1847
rect 3002 1327 3010 1332
rect 3040 1707 3056 1902
rect 3045 1702 3050 1707
rect 3055 1702 3056 1707
rect 3040 1507 3056 1702
rect 3045 1502 3050 1507
rect 3055 1502 3056 1507
rect 3040 1307 3056 1502
rect 3045 1302 3050 1307
rect 3055 1302 3056 1307
rect 3040 1107 3056 1302
rect 3045 1102 3050 1107
rect 3055 1102 3056 1107
rect 3040 907 3056 1102
rect 3045 902 3050 907
rect 3055 902 3056 907
rect 3040 707 3056 902
rect 3045 702 3050 707
rect 3055 702 3056 707
rect 3040 507 3056 702
rect 3045 502 3050 507
rect 3055 502 3056 507
rect 2541 202 2546 207
rect 2551 202 2552 207
rect 2536 7 2552 202
rect 2765 22 2770 317
rect 3040 307 3056 502
rect 3045 302 3050 307
rect 3055 302 3056 307
rect 3040 107 3056 302
rect 3045 102 3050 107
rect 3055 102 3056 107
rect 2541 2 2546 7
rect 2551 2 2552 7
rect 2536 -30 2552 2
rect 3040 -30 3056 102
rect 3325 72 3330 1477
rect 3357 72 3362 1557
rect 3437 382 3442 3257
rect 3453 2332 3458 3237
rect 3469 1552 3474 2357
rect 3485 1582 3490 2157
rect 3501 1612 3506 3287
rect 3485 82 3490 1337
rect 3517 992 3522 1687
use BUFX4  BUFX4_54
timestamp 1696145522
transform 1 0 36 0 1 105
box -2 -3 34 103
use BUFX4  BUFX4_44
timestamp 1696145522
transform 1 0 4 0 1 105
box -2 -3 34 103
use BUFX4  BUFX4_48
timestamp 1696145522
transform 1 0 36 0 -1 105
box -2 -3 34 103
use BUFX4  BUFX4_49
timestamp 1696145522
transform 1 0 4 0 -1 105
box -2 -3 34 103
use BUFX4  BUFX4_53
timestamp 1696145522
transform 1 0 68 0 1 105
box -2 -3 34 103
use BUFX4  BUFX4_52
timestamp 1696145522
transform 1 0 68 0 -1 105
box -2 -3 34 103
use BUFX4  BUFX4_187
timestamp 1696145522
transform -1 0 132 0 1 105
box -2 -3 34 103
use BUFX4  BUFX4_47
timestamp 1696145522
transform 1 0 100 0 -1 105
box -2 -3 34 103
use BUFX4  BUFX4_188
timestamp 1696145522
transform 1 0 132 0 1 105
box -2 -3 34 103
use BUFX4  BUFX4_193
timestamp 1696145522
transform 1 0 132 0 -1 105
box -2 -3 34 103
use BUFX4  BUFX4_190
timestamp 1696145522
transform 1 0 164 0 1 105
box -2 -3 34 103
use BUFX2  BUFX2_1
timestamp 1696145522
transform -1 0 188 0 -1 105
box -2 -3 26 103
use BUFX4  BUFX4_189
timestamp 1696145522
transform 1 0 196 0 1 105
box -2 -3 34 103
use BUFX4  BUFX4_130
timestamp 1696145522
transform 1 0 212 0 -1 105
box -2 -3 34 103
use BUFX2  BUFX2_2
timestamp 1696145522
transform 1 0 188 0 -1 105
box -2 -3 26 103
use BUFX4  BUFX4_55
timestamp 1696145522
transform 1 0 228 0 1 105
box -2 -3 34 103
use BUFX4  BUFX4_46
timestamp 1696145522
transform 1 0 244 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_220
timestamp 1696145522
transform 1 0 292 0 1 105
box -2 -3 26 103
use BUFX4  BUFX4_45
timestamp 1696145522
transform 1 0 260 0 1 105
box -2 -3 34 103
use BUFX4  BUFX4_35
timestamp 1696145522
transform 1 0 276 0 -1 105
box -2 -3 34 103
use BUFX4  BUFX4_76
timestamp 1696145522
transform 1 0 316 0 1 105
box -2 -3 34 103
use BUFX4  BUFX4_74
timestamp 1696145522
transform 1 0 308 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_120
timestamp 1696145522
transform 1 0 348 0 1 105
box -2 -3 34 103
use INVX1  INVX1_68
timestamp 1696145522
transform -1 0 380 0 -1 105
box -2 -3 18 103
use NAND2X1  NAND2X1_107
timestamp 1696145522
transform 1 0 340 0 -1 105
box -2 -3 26 103
use INVX8  INVX8_1
timestamp 1696145522
transform -1 0 420 0 1 105
box -2 -3 42 103
use NAND2X1  NAND2X1_238
timestamp 1696145522
transform 1 0 412 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_117
timestamp 1696145522
transform 1 0 380 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_164
timestamp 1696145522
transform -1 0 476 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_207
timestamp 1696145522
transform -1 0 452 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_224
timestamp 1696145522
transform 1 0 460 0 -1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_161
timestamp 1696145522
transform 1 0 436 0 -1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_103
timestamp 1696145522
transform 1 0 524 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_191
timestamp 1696145522
transform -1 0 524 0 1 105
box -2 -3 34 103
use FILL  FILL_1_0_1
timestamp 1696145522
transform -1 0 492 0 1 105
box -2 -3 10 103
use FILL  FILL_1_0_0
timestamp 1696145522
transform -1 0 484 0 1 105
box -2 -3 10 103
use MUX2X1  MUX2X1_12
timestamp 1696145522
transform -1 0 548 0 -1 105
box -2 -3 50 103
use FILL  FILL_0_0_1
timestamp 1696145522
transform -1 0 500 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_0_0
timestamp 1696145522
transform -1 0 492 0 -1 105
box -2 -3 10 103
use OAI21X1  OAI21X1_190
timestamp 1696145522
transform -1 0 628 0 1 105
box -2 -3 34 103
use MUX2X1  MUX2X1_4
timestamp 1696145522
transform 1 0 548 0 1 105
box -2 -3 50 103
use NAND2X1  NAND2X1_242
timestamp 1696145522
transform 1 0 580 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_211
timestamp 1696145522
transform 1 0 548 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_114
timestamp 1696145522
transform 1 0 628 0 1 105
box -2 -3 34 103
use MUX2X1  MUX2X1_11
timestamp 1696145522
transform -1 0 676 0 -1 105
box -2 -3 50 103
use NAND2X1  NAND2X1_104
timestamp 1696145522
transform 1 0 604 0 -1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_560
timestamp 1696145522
transform 1 0 684 0 1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_158
timestamp 1696145522
transform 1 0 660 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_57
timestamp 1696145522
transform -1 0 732 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_106
timestamp 1696145522
transform 1 0 676 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_682
timestamp 1696145522
transform -1 0 740 0 1 105
box -2 -3 34 103
use MUX2X1  MUX2X1_3
timestamp 1696145522
transform -1 0 820 0 1 105
box -2 -3 50 103
use INVX1  INVX1_44
timestamp 1696145522
transform -1 0 772 0 1 105
box -2 -3 18 103
use INVX1  INVX1_286
timestamp 1696145522
transform 1 0 740 0 1 105
box -2 -3 18 103
use NAND2X1  NAND2X1_562
timestamp 1696145522
transform 1 0 764 0 -1 105
box -2 -3 26 103
use BUFX4  BUFX4_66
timestamp 1696145522
transform 1 0 732 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_579
timestamp 1696145522
transform -1 0 844 0 1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_102
timestamp 1696145522
transform 1 0 820 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_689
timestamp 1696145522
transform -1 0 820 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_241
timestamp 1696145522
transform -1 0 900 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_53
timestamp 1696145522
transform -1 0 876 0 1 105
box -2 -3 34 103
use MUX2X1  MUX2X1_1
timestamp 1696145522
transform 1 0 868 0 -1 105
box -2 -3 50 103
use NAND2X1  NAND2X1_100
timestamp 1696145522
transform 1 0 844 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_51
timestamp 1696145522
transform -1 0 932 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_155
timestamp 1696145522
transform 1 0 956 0 1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_76
timestamp 1696145522
transform 1 0 932 0 1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_162
timestamp 1696145522
transform 1 0 964 0 -1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_297
timestamp 1696145522
transform -1 0 964 0 -1 105
box -2 -3 34 103
use INVX2  INVX2_58
timestamp 1696145522
transform -1 0 932 0 -1 105
box -2 -3 18 103
use XOR2X1  XOR2X1_3
timestamp 1696145522
transform 1 0 996 0 1 105
box -2 -3 58 103
use FILL  FILL_1_1_1
timestamp 1696145522
transform 1 0 988 0 1 105
box -2 -3 10 103
use FILL  FILL_1_1_0
timestamp 1696145522
transform 1 0 980 0 1 105
box -2 -3 10 103
use OAI21X1  OAI21X1_118
timestamp 1696145522
transform -1 0 1036 0 -1 105
box -2 -3 34 103
use FILL  FILL_0_1_1
timestamp 1696145522
transform -1 0 1004 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_1_0
timestamp 1696145522
transform -1 0 996 0 -1 105
box -2 -3 10 103
use MUX2X1  MUX2X1_89
timestamp 1696145522
transform 1 0 1052 0 1 105
box -2 -3 50 103
use OAI21X1  OAI21X1_116
timestamp 1696145522
transform -1 0 1092 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_160
timestamp 1696145522
transform 1 0 1036 0 -1 105
box -2 -3 26 103
use MUX2X1  MUX2X1_84
timestamp 1696145522
transform 1 0 1148 0 1 105
box -2 -3 50 103
use MUX2X1  MUX2X1_91
timestamp 1696145522
transform 1 0 1100 0 1 105
box -2 -3 50 103
use XNOR2X1  XNOR2X1_16
timestamp 1696145522
transform 1 0 1124 0 -1 105
box -2 -3 58 103
use INVX2  INVX2_13
timestamp 1696145522
transform 1 0 1108 0 -1 105
box -2 -3 18 103
use INVX2  INVX2_20
timestamp 1696145522
transform -1 0 1108 0 -1 105
box -2 -3 18 103
use INVX2  INVX2_12
timestamp 1696145522
transform 1 0 1196 0 1 105
box -2 -3 18 103
use NOR2X1  NOR2X1_112
timestamp 1696145522
transform -1 0 1220 0 -1 105
box -2 -3 26 103
use INVX1  INVX1_79
timestamp 1696145522
transform 1 0 1180 0 -1 105
box -2 -3 18 103
use MUX2X1  MUX2X1_82
timestamp 1696145522
transform -1 0 1300 0 1 105
box -2 -3 50 103
use NAND2X1  NAND2X1_68
timestamp 1696145522
transform -1 0 1252 0 1 105
box -2 -3 26 103
use INVX1  INVX1_29
timestamp 1696145522
transform 1 0 1212 0 1 105
box -2 -3 18 103
use OAI21X1  OAI21X1_642
timestamp 1696145522
transform 1 0 1244 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_194
timestamp 1696145522
transform 1 0 1220 0 -1 105
box -2 -3 26 103
use MUX2X1  MUX2X1_85
timestamp 1696145522
transform -1 0 1348 0 1 105
box -2 -3 50 103
use XNOR2X1  XNOR2X1_17
timestamp 1696145522
transform 1 0 1292 0 -1 105
box -2 -3 58 103
use INVX1  INVX1_279
timestamp 1696145522
transform -1 0 1292 0 -1 105
box -2 -3 18 103
use NOR2X1  NOR2X1_54
timestamp 1696145522
transform 1 0 1380 0 1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_22
timestamp 1696145522
transform 1 0 1348 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_69
timestamp 1696145522
transform 1 0 1380 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_156
timestamp 1696145522
transform 1 0 1348 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_28
timestamp 1696145522
transform 1 0 1444 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_67
timestamp 1696145522
transform -1 0 1444 0 1 105
box -2 -3 26 103
use INVX2  INVX2_9
timestamp 1696145522
transform 1 0 1404 0 1 105
box -2 -3 18 103
use OAI21X1  OAI21X1_713
timestamp 1696145522
transform 1 0 1436 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_643
timestamp 1696145522
transform 1 0 1404 0 -1 105
box -2 -3 34 103
use FILL  FILL_1_2_0
timestamp 1696145522
transform 1 0 1508 0 1 105
box -2 -3 10 103
use AOI21X1  AOI21X1_277
timestamp 1696145522
transform 1 0 1476 0 1 105
box -2 -3 34 103
use INVX2  INVX2_26
timestamp 1696145522
transform -1 0 1516 0 -1 105
box -2 -3 18 103
use AOI21X1  AOI21X1_304
timestamp 1696145522
transform 1 0 1468 0 -1 105
box -2 -3 34 103
use AOI21X1  AOI21X1_312
timestamp 1696145522
transform 1 0 1556 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_743
timestamp 1696145522
transform 1 0 1524 0 1 105
box -2 -3 34 103
use FILL  FILL_1_2_1
timestamp 1696145522
transform 1 0 1516 0 1 105
box -2 -3 10 103
use XNOR2X1  XNOR2X1_18
timestamp 1696145522
transform -1 0 1620 0 -1 105
box -2 -3 58 103
use AOI21X1  AOI21X1_306
timestamp 1696145522
transform 1 0 1532 0 -1 105
box -2 -3 34 103
use FILL  FILL_0_2_1
timestamp 1696145522
transform 1 0 1524 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_2_0
timestamp 1696145522
transform 1 0 1516 0 -1 105
box -2 -3 10 103
use NOR2X1  NOR2X1_107
timestamp 1696145522
transform -1 0 1644 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_744
timestamp 1696145522
transform -1 0 1620 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_58
timestamp 1696145522
transform -1 0 1644 0 -1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_51
timestamp 1696145522
transform -1 0 1708 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_729
timestamp 1696145522
transform -1 0 1676 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_20
timestamp 1696145522
transform 1 0 1676 0 -1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_25
timestamp 1696145522
transform 1 0 1644 0 -1 105
box -2 -3 34 103
use AND2X2  AND2X2_46
timestamp 1696145522
transform 1 0 1732 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_410
timestamp 1696145522
transform 1 0 1708 0 1 105
box -2 -3 26 103
use INVX1  INVX1_13
timestamp 1696145522
transform 1 0 1740 0 -1 105
box -2 -3 18 103
use NOR2X1  NOR2X1_25
timestamp 1696145522
transform -1 0 1740 0 -1 105
box -2 -3 26 103
use INVX1  INVX1_12
timestamp 1696145522
transform 1 0 1700 0 -1 105
box -2 -3 18 103
use XNOR2X1  XNOR2X1_19
timestamp 1696145522
transform 1 0 1764 0 1 105
box -2 -3 58 103
use INVX1  INVX1_281
timestamp 1696145522
transform 1 0 1804 0 -1 105
box -2 -3 18 103
use NAND2X1  NAND2X1_22
timestamp 1696145522
transform 1 0 1780 0 -1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_21
timestamp 1696145522
transform -1 0 1780 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_774
timestamp 1696145522
transform 1 0 1852 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_787
timestamp 1696145522
transform 1 0 1820 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_10
timestamp 1696145522
transform 1 0 1844 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_23
timestamp 1696145522
transform -1 0 1844 0 -1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_26
timestamp 1696145522
transform 1 0 1924 0 1 105
box -2 -3 26 103
use INVX1  INVX1_14
timestamp 1696145522
transform 1 0 1908 0 1 105
box -2 -3 18 103
use NAND2X1  NAND2X1_21
timestamp 1696145522
transform 1 0 1884 0 1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_279
timestamp 1696145522
transform -1 0 1956 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_159
timestamp 1696145522
transform -1 0 1924 0 -1 105
box -2 -3 34 103
use INVX1  INVX1_81
timestamp 1696145522
transform 1 0 1876 0 -1 105
box -2 -3 18 103
use XOR2X1  XOR2X1_5
timestamp 1696145522
transform -1 0 2004 0 1 105
box -2 -3 58 103
use NOR2X1  NOR2X1_114
timestamp 1696145522
transform -1 0 2012 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_783
timestamp 1696145522
transform -1 0 1988 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_158
timestamp 1696145522
transform -1 0 2076 0 1 105
box -2 -3 34 103
use FILL  FILL_1_3_1
timestamp 1696145522
transform -1 0 2044 0 1 105
box -2 -3 10 103
use FILL  FILL_1_3_0
timestamp 1696145522
transform -1 0 2036 0 1 105
box -2 -3 10 103
use NAND2X1  NAND2X1_71
timestamp 1696145522
transform 1 0 2004 0 1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_52
timestamp 1696145522
transform -1 0 2060 0 -1 105
box -2 -3 34 103
use FILL  FILL_0_3_1
timestamp 1696145522
transform -1 0 2028 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_3_0
timestamp 1696145522
transform -1 0 2020 0 -1 105
box -2 -3 10 103
use OAI21X1  OAI21X1_644
timestamp 1696145522
transform 1 0 2108 0 1 105
box -2 -3 34 103
use AOI21X1  AOI21X1_278
timestamp 1696145522
transform 1 0 2076 0 1 105
box -2 -3 34 103
use INVX2  INVX2_24
timestamp 1696145522
transform -1 0 2132 0 -1 105
box -2 -3 18 103
use XNOR2X1  XNOR2X1_40
timestamp 1696145522
transform 1 0 2060 0 -1 105
box -2 -3 58 103
use AOI21X1  AOI21X1_26
timestamp 1696145522
transform -1 0 2204 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_29
timestamp 1696145522
transform -1 0 2172 0 1 105
box -2 -3 34 103
use XNOR2X1  XNOR2X1_9
timestamp 1696145522
transform 1 0 2156 0 -1 105
box -2 -3 58 103
use BUFX2  BUFX2_7
timestamp 1696145522
transform -1 0 2156 0 -1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_56
timestamp 1696145522
transform 1 0 2204 0 1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_62
timestamp 1696145522
transform 1 0 2212 0 -1 105
box -2 -3 26 103
use OR2X2  OR2X2_3
timestamp 1696145522
transform 1 0 2228 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_539
timestamp 1696145522
transform 1 0 2236 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_160
timestamp 1696145522
transform -1 0 2292 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_38
timestamp 1696145522
transform -1 0 2308 0 -1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_64
timestamp 1696145522
transform -1 0 2284 0 -1 105
box -2 -3 26 103
use AND2X2  AND2X2_47
timestamp 1696145522
transform 1 0 2292 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_35
timestamp 1696145522
transform 1 0 2308 0 -1 105
box -2 -3 26 103
use NAND3X1  NAND3X1_52
timestamp 1696145522
transform 1 0 2356 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_645
timestamp 1696145522
transform 1 0 2324 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_32
timestamp 1696145522
transform -1 0 2380 0 -1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_41
timestamp 1696145522
transform 1 0 2332 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_798
timestamp 1696145522
transform -1 0 2420 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_79
timestamp 1696145522
transform -1 0 2436 0 -1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_27
timestamp 1696145522
transform 1 0 2380 0 -1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_33
timestamp 1696145522
transform -1 0 2484 0 1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_202
timestamp 1696145522
transform 1 0 2436 0 1 105
box -2 -3 26 103
use INVX1  INVX1_20
timestamp 1696145522
transform 1 0 2420 0 1 105
box -2 -3 18 103
use XNOR2X1  XNOR2X1_8
timestamp 1696145522
transform -1 0 2532 0 -1 105
box -2 -3 58 103
use INVX2  INVX2_25
timestamp 1696145522
transform -1 0 2476 0 -1 105
box -2 -3 18 103
use NOR2X1  NOR2X1_61
timestamp 1696145522
transform -1 0 2460 0 -1 105
box -2 -3 26 103
use XNOR2X1  XNOR2X1_5
timestamp 1696145522
transform 1 0 2532 0 1 105
box -2 -3 58 103
use FILL  FILL_1_4_1
timestamp 1696145522
transform 1 0 2524 0 1 105
box -2 -3 10 103
use FILL  FILL_1_4_0
timestamp 1696145522
transform 1 0 2516 0 1 105
box -2 -3 10 103
use INVX1  INVX1_21
timestamp 1696145522
transform 1 0 2500 0 1 105
box -2 -3 18 103
use INVX1  INVX1_278
timestamp 1696145522
transform 1 0 2484 0 1 105
box -2 -3 18 103
use FILL  FILL_0_4_0
timestamp 1696145522
transform -1 0 2540 0 -1 105
box -2 -3 10 103
use NOR2X1  NOR2X1_36
timestamp 1696145522
transform 1 0 2588 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_161
timestamp 1696145522
transform 1 0 2596 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_201
timestamp 1696145522
transform 1 0 2572 0 -1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_117
timestamp 1696145522
transform -1 0 2572 0 -1 105
box -2 -3 26 103
use FILL  FILL_0_4_1
timestamp 1696145522
transform -1 0 2548 0 -1 105
box -2 -3 10 103
use NAND2X1  NAND2X1_36
timestamp 1696145522
transform 1 0 2652 0 1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_34
timestamp 1696145522
transform -1 0 2652 0 1 105
box -2 -3 26 103
use INVX1  INVX1_18
timestamp 1696145522
transform 1 0 2612 0 1 105
box -2 -3 18 103
use OAI21X1  OAI21X1_639
timestamp 1696145522
transform -1 0 2660 0 -1 105
box -2 -3 34 103
use XNOR2X1  XNOR2X1_4
timestamp 1696145522
transform -1 0 2732 0 1 105
box -2 -3 58 103
use AND2X2  AND2X2_10
timestamp 1696145522
transform -1 0 2724 0 -1 105
box -2 -3 34 103
use AOI21X1  AOI21X1_55
timestamp 1696145522
transform 1 0 2660 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_806
timestamp 1696145522
transform -1 0 2788 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_65
timestamp 1696145522
transform 1 0 2732 0 1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_78
timestamp 1696145522
transform 1 0 2756 0 -1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_343
timestamp 1696145522
transform 1 0 2724 0 -1 105
box -2 -3 34 103
use AOI21X1  AOI21X1_29
timestamp 1696145522
transform -1 0 2844 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_77
timestamp 1696145522
transform -1 0 2812 0 1 105
box -2 -3 26 103
use XNOR2X1  XNOR2X1_7
timestamp 1696145522
transform -1 0 2860 0 -1 105
box -2 -3 58 103
use NOR2X1  NOR2X1_60
timestamp 1696145522
transform -1 0 2804 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_818
timestamp 1696145522
transform 1 0 2876 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_641
timestamp 1696145522
transform -1 0 2876 0 1 105
box -2 -3 34 103
use XNOR2X1  XNOR2X1_22
timestamp 1696145522
transform 1 0 2860 0 -1 105
box -2 -3 58 103
use NAND2X1  NAND2X1_75
timestamp 1696145522
transform 1 0 2956 0 1 105
box -2 -3 26 103
use INVX2  INVX2_15
timestamp 1696145522
transform -1 0 2956 0 1 105
box -2 -3 18 103
use OAI21X1  OAI21X1_32
timestamp 1696145522
transform 1 0 2908 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_164
timestamp 1696145522
transform -1 0 2980 0 -1 105
box -2 -3 34 103
use AOI21X1  AOI21X1_53
timestamp 1696145522
transform 1 0 2916 0 -1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_640
timestamp 1696145522
transform 1 0 3020 0 1 105
box -2 -3 34 103
use AOI22X1  AOI22X1_29
timestamp 1696145522
transform 1 0 2980 0 1 105
box -2 -3 42 103
use XOR2X1  XOR2X1_8
timestamp 1696145522
transform 1 0 2980 0 -1 105
box -2 -3 58 103
use NAND2X1  NAND2X1_76
timestamp 1696145522
transform -1 0 3092 0 1 105
box -2 -3 26 103
use FILL  FILL_1_5_1
timestamp 1696145522
transform -1 0 3068 0 1 105
box -2 -3 10 103
use FILL  FILL_1_5_0
timestamp 1696145522
transform -1 0 3060 0 1 105
box -2 -3 10 103
use XOR2X1  XOR2X1_6
timestamp 1696145522
transform 1 0 3076 0 -1 105
box -2 -3 58 103
use FILL  FILL_0_5_1
timestamp 1696145522
transform 1 0 3068 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_5_0
timestamp 1696145522
transform 1 0 3060 0 -1 105
box -2 -3 10 103
use NOR2X1  NOR2X1_116
timestamp 1696145522
transform -1 0 3060 0 -1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_31
timestamp 1696145522
transform 1 0 3124 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_30
timestamp 1696145522
transform 1 0 3092 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_59
timestamp 1696145522
transform -1 0 3156 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_31
timestamp 1696145522
transform 1 0 3172 0 1 105
box -2 -3 34 103
use INVX1  INVX1_82
timestamp 1696145522
transform 1 0 3156 0 1 105
box -2 -3 18 103
use XNOR2X1  XNOR2X1_6
timestamp 1696145522
transform 1 0 3156 0 -1 105
box -2 -3 58 103
use AOI21X1  AOI21X1_353
timestamp 1696145522
transform 1 0 3244 0 1 105
box -2 -3 34 103
use INVX1  INVX1_314
timestamp 1696145522
transform 1 0 3228 0 1 105
box -2 -3 18 103
use NAND2X1  NAND2X1_200
timestamp 1696145522
transform -1 0 3228 0 1 105
box -2 -3 26 103
use XNOR2X1  XNOR2X1_44
timestamp 1696145522
transform -1 0 3292 0 -1 105
box -2 -3 58 103
use NAND2X1  NAND2X1_64
timestamp 1696145522
transform -1 0 3236 0 -1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_28
timestamp 1696145522
transform -1 0 3380 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_74
timestamp 1696145522
transform 1 0 3324 0 1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_54
timestamp 1696145522
transform 1 0 3292 0 1 105
box -2 -3 34 103
use INVX1  INVX1_84
timestamp 1696145522
transform 1 0 3276 0 1 105
box -2 -3 18 103
use INVX4  INVX4_4
timestamp 1696145522
transform -1 0 3372 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_902
timestamp 1696145522
transform -1 0 3348 0 -1 105
box -2 -3 34 103
use BUFX2  BUFX2_24
timestamp 1696145522
transform 1 0 3292 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_162
timestamp 1696145522
transform -1 0 3460 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_638
timestamp 1696145522
transform -1 0 3428 0 1 105
box -2 -3 34 103
use INVX1  INVX1_83
timestamp 1696145522
transform 1 0 3380 0 1 105
box -2 -3 18 103
use DFFSR  DFFSR_1
timestamp 1696145522
transform -1 0 3548 0 -1 105
box -2 -3 178 103
use FILL  FILL_1_1
timestamp 1696145522
transform -1 0 3556 0 -1 105
box -2 -3 10 103
use FILL  FILL_1_2
timestamp 1696145522
transform -1 0 3564 0 -1 105
box -2 -3 10 103
use NOR2X1  NOR2X1_118
timestamp 1696145522
transform 1 0 3460 0 1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_63
timestamp 1696145522
transform 1 0 3484 0 1 105
box -2 -3 26 103
use INVX2  INVX2_27
timestamp 1696145522
transform 1 0 3508 0 1 105
box -2 -3 18 103
use AOI21X1  AOI21X1_58
timestamp 1696145522
transform -1 0 3556 0 1 105
box -2 -3 34 103
use FILL  FILL_2_1
timestamp 1696145522
transform 1 0 3556 0 1 105
box -2 -3 10 103
use BUFX4  BUFX4_51
timestamp 1696145522
transform 1 0 4 0 -1 305
box -2 -3 34 103
use BUFX4  BUFX4_43
timestamp 1696145522
transform 1 0 36 0 -1 305
box -2 -3 34 103
use BUFX4  BUFX4_50
timestamp 1696145522
transform 1 0 68 0 -1 305
box -2 -3 34 103
use BUFX4  BUFX4_194
timestamp 1696145522
transform -1 0 132 0 -1 305
box -2 -3 34 103
use BUFX4  BUFX4_191
timestamp 1696145522
transform 1 0 132 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_222
timestamp 1696145522
transform 1 0 164 0 -1 305
box -2 -3 26 103
use BUFX4  BUFX4_196
timestamp 1696145522
transform 1 0 188 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_105
timestamp 1696145522
transform 1 0 220 0 -1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_221
timestamp 1696145522
transform 1 0 244 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_187
timestamp 1696145522
transform 1 0 268 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_308
timestamp 1696145522
transform -1 0 324 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_58
timestamp 1696145522
transform 1 0 324 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_277
timestamp 1696145522
transform -1 0 380 0 -1 305
box -2 -3 26 103
use INVX1  INVX1_67
timestamp 1696145522
transform -1 0 396 0 -1 305
box -2 -3 18 103
use NAND2X1  NAND2X1_302
timestamp 1696145522
transform -1 0 420 0 -1 305
box -2 -3 26 103
use MUX2X1  MUX2X1_35
timestamp 1696145522
transform -1 0 468 0 -1 305
box -2 -3 50 103
use NAND2X1  NAND2X1_225
timestamp 1696145522
transform 1 0 468 0 -1 305
box -2 -3 26 103
use FILL  FILL_2_0_0
timestamp 1696145522
transform 1 0 492 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_0_1
timestamp 1696145522
transform 1 0 500 0 -1 305
box -2 -3 10 103
use OAI21X1  OAI21X1_290
timestamp 1696145522
transform 1 0 508 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_54
timestamp 1696145522
transform -1 0 572 0 -1 305
box -2 -3 34 103
use INVX1  INVX1_90
timestamp 1696145522
transform -1 0 588 0 -1 305
box -2 -3 18 103
use NAND2X1  NAND2X1_223
timestamp 1696145522
transform 1 0 588 0 -1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_85
timestamp 1696145522
transform 1 0 612 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_55
timestamp 1696145522
transform -1 0 668 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_561
timestamp 1696145522
transform 1 0 668 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_684
timestamp 1696145522
transform -1 0 724 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_683
timestamp 1696145522
transform -1 0 756 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_577
timestamp 1696145522
transform -1 0 780 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_685
timestamp 1696145522
transform -1 0 812 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_719
timestamp 1696145522
transform 1 0 812 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_243
timestamp 1696145522
transform -1 0 868 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_210
timestamp 1696145522
transform -1 0 900 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_690
timestamp 1696145522
transform -1 0 932 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_156
timestamp 1696145522
transform 1 0 932 0 -1 305
box -2 -3 26 103
use INVX1  INVX1_65
timestamp 1696145522
transform -1 0 972 0 -1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_111
timestamp 1696145522
transform -1 0 1004 0 -1 305
box -2 -3 34 103
use FILL  FILL_2_1_0
timestamp 1696145522
transform 1 0 1004 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_1_1
timestamp 1696145522
transform 1 0 1012 0 -1 305
box -2 -3 10 103
use NOR2X1  NOR2X1_432
timestamp 1696145522
transform 1 0 1020 0 -1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_298
timestamp 1696145522
transform 1 0 1044 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_692
timestamp 1696145522
transform -1 0 1108 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_52
timestamp 1696145522
transform 1 0 1108 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_691
timestamp 1696145522
transform -1 0 1172 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_101
timestamp 1696145522
transform 1 0 1172 0 -1 305
box -2 -3 26 103
use MUX2X1  MUX2X1_92
timestamp 1696145522
transform -1 0 1244 0 -1 305
box -2 -3 50 103
use OAI21X1  OAI21X1_119
timestamp 1696145522
transform -1 0 1276 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_157
timestamp 1696145522
transform 1 0 1276 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_113
timestamp 1696145522
transform -1 0 1332 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_20
timestamp 1696145522
transform 1 0 1332 0 -1 305
box -2 -3 26 103
use NOR2X1  NOR2X1_408
timestamp 1696145522
transform -1 0 1380 0 -1 305
box -2 -3 26 103
use NOR2X1  NOR2X1_15
timestamp 1696145522
transform 1 0 1380 0 -1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_48
timestamp 1696145522
transform 1 0 1404 0 -1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_18
timestamp 1696145522
transform 1 0 1436 0 -1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_23
timestamp 1696145522
transform -1 0 1492 0 -1 305
box -2 -3 34 103
use INVX1  INVX1_280
timestamp 1696145522
transform 1 0 1492 0 -1 305
box -2 -3 18 103
use FILL  FILL_2_2_0
timestamp 1696145522
transform 1 0 1508 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_2_1
timestamp 1696145522
transform 1 0 1516 0 -1 305
box -2 -3 10 103
use NOR2X1  NOR2X1_19
timestamp 1696145522
transform 1 0 1524 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_8
timestamp 1696145522
transform 1 0 1548 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_199
timestamp 1696145522
transform 1 0 1580 0 -1 305
box -2 -3 26 103
use INVX1  INVX1_80
timestamp 1696145522
transform 1 0 1604 0 -1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_157
timestamp 1696145522
transform -1 0 1652 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_152
timestamp 1696145522
transform -1 0 1684 0 -1 305
box -2 -3 34 103
use INVX4  INVX4_7
timestamp 1696145522
transform 1 0 1684 0 -1 305
box -2 -3 26 103
use NOR2X1  NOR2X1_113
timestamp 1696145522
transform 1 0 1708 0 -1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_307
timestamp 1696145522
transform 1 0 1732 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_9
timestamp 1696145522
transform 1 0 1764 0 -1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_49
timestamp 1696145522
transform 1 0 1796 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_788
timestamp 1696145522
transform -1 0 1860 0 -1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_316
timestamp 1696145522
transform -1 0 1892 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_752
timestamp 1696145522
transform -1 0 1924 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_26
timestamp 1696145522
transform 1 0 1924 0 -1 305
box -2 -3 26 103
use INVX2  INVX2_92
timestamp 1696145522
transform 1 0 1948 0 -1 305
box -2 -3 18 103
use INVX1  INVX1_298
timestamp 1696145522
transform 1 0 1964 0 -1 305
box -2 -3 18 103
use NAND3X1  NAND3X1_4
timestamp 1696145522
transform -1 0 2012 0 -1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_108
timestamp 1696145522
transform 1 0 2012 0 -1 305
box -2 -3 26 103
use FILL  FILL_2_3_0
timestamp 1696145522
transform -1 0 2044 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_3_1
timestamp 1696145522
transform -1 0 2052 0 -1 305
box -2 -3 10 103
use OAI21X1  OAI21X1_758
timestamp 1696145522
transform -1 0 2084 0 -1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_317
timestamp 1696145522
transform -1 0 2116 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_757
timestamp 1696145522
transform -1 0 2148 0 -1 305
box -2 -3 34 103
use XNOR2X1  XNOR2X1_20
timestamp 1696145522
transform -1 0 2204 0 -1 305
box -2 -3 58 103
use NAND2X1  NAND2X1_72
timestamp 1696145522
transform -1 0 2228 0 -1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_759
timestamp 1696145522
transform 1 0 2228 0 -1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_318
timestamp 1696145522
transform 1 0 2260 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_772
timestamp 1696145522
transform 1 0 2292 0 -1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_8
timestamp 1696145522
transform -1 0 2356 0 -1 305
box -2 -3 34 103
use BUFX2  BUFX2_6
timestamp 1696145522
transform 1 0 2356 0 -1 305
box -2 -3 26 103
use NOR2X1  NOR2X1_448
timestamp 1696145522
transform 1 0 2380 0 -1 305
box -2 -3 26 103
use BUFX2  BUFX2_8
timestamp 1696145522
transform 1 0 2404 0 -1 305
box -2 -3 26 103
use INVX1  INVX1_302
timestamp 1696145522
transform -1 0 2444 0 -1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_773
timestamp 1696145522
transform 1 0 2444 0 -1 305
box -2 -3 34 103
use AOI22X1  AOI22X1_36
timestamp 1696145522
transform -1 0 2516 0 -1 305
box -2 -3 42 103
use AOI21X1  AOI21X1_328
timestamp 1696145522
transform -1 0 2548 0 -1 305
box -2 -3 34 103
use FILL  FILL_2_4_0
timestamp 1696145522
transform 1 0 2548 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_4_1
timestamp 1696145522
transform 1 0 2556 0 -1 305
box -2 -3 10 103
use OAI21X1  OAI21X1_838
timestamp 1696145522
transform 1 0 2564 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_837
timestamp 1696145522
transform -1 0 2628 0 -1 305
box -2 -3 34 103
use INVX2  INVX2_21
timestamp 1696145522
transform -1 0 2644 0 -1 305
box -2 -3 18 103
use NAND2X1  NAND2X1_37
timestamp 1696145522
transform 1 0 2644 0 -1 305
box -2 -3 26 103
use INVX1  INVX1_19
timestamp 1696145522
transform -1 0 2684 0 -1 305
box -2 -3 18 103
use NOR2X1  NOR2X1_37
timestamp 1696145522
transform -1 0 2708 0 -1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_38
timestamp 1696145522
transform 1 0 2708 0 -1 305
box -2 -3 26 103
use XNOR2X1  XNOR2X1_41
timestamp 1696145522
transform -1 0 2788 0 -1 305
box -2 -3 58 103
use AOI21X1  AOI21X1_345
timestamp 1696145522
transform 1 0 2788 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_845
timestamp 1696145522
transform -1 0 2852 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_39
timestamp 1696145522
transform 1 0 2852 0 -1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_40
timestamp 1696145522
transform 1 0 2876 0 -1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_344
timestamp 1696145522
transform 1 0 2900 0 -1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_834
timestamp 1696145522
transform 1 0 2932 0 -1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_27
timestamp 1696145522
transform 1 0 2964 0 -1 305
box -2 -3 26 103
use AND2X2  AND2X2_48
timestamp 1696145522
transform 1 0 2988 0 -1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_115
timestamp 1696145522
transform -1 0 3044 0 -1 305
box -2 -3 26 103
use FILL  FILL_2_5_0
timestamp 1696145522
transform -1 0 3052 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_5_1
timestamp 1696145522
transform -1 0 3060 0 -1 305
box -2 -3 10 103
use NOR2X1  NOR2X1_39
timestamp 1696145522
transform -1 0 3084 0 -1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_43
timestamp 1696145522
transform 1 0 3084 0 -1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_28
timestamp 1696145522
transform 1 0 3108 0 -1 305
box -2 -3 26 103
use INVX1  INVX1_15
timestamp 1696145522
transform -1 0 3148 0 -1 305
box -2 -3 18 103
use NAND2X1  NAND2X1_29
timestamp 1696145522
transform -1 0 3172 0 -1 305
box -2 -3 26 103
use INVX1  INVX1_30
timestamp 1696145522
transform -1 0 3188 0 -1 305
box -2 -3 18 103
use AOI21X1  AOI21X1_30
timestamp 1696145522
transform -1 0 3220 0 -1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_30
timestamp 1696145522
transform -1 0 3244 0 -1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_280
timestamp 1696145522
transform 1 0 3244 0 -1 305
box -2 -3 34 103
use INVX1  INVX1_85
timestamp 1696145522
transform 1 0 3276 0 -1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_163
timestamp 1696145522
transform 1 0 3292 0 -1 305
box -2 -3 34 103
use XNOR2X1  XNOR2X1_23
timestamp 1696145522
transform -1 0 3380 0 -1 305
box -2 -3 58 103
use OAI21X1  OAI21X1_16
timestamp 1696145522
transform -1 0 3412 0 -1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_30
timestamp 1696145522
transform 1 0 3412 0 -1 305
box -2 -3 26 103
use INVX2  INVX2_23
timestamp 1696145522
transform 1 0 3436 0 -1 305
box -2 -3 18 103
use NAND2X1  NAND2X1_203
timestamp 1696145522
transform -1 0 3476 0 -1 305
box -2 -3 26 103
use NOR2X1  NOR2X1_31
timestamp 1696145522
transform 1 0 3476 0 -1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_42
timestamp 1696145522
transform -1 0 3524 0 -1 305
box -2 -3 26 103
use NOR2X1  NOR2X1_34
timestamp 1696145522
transform 1 0 3524 0 -1 305
box -2 -3 26 103
use FILL  FILL_3_1
timestamp 1696145522
transform -1 0 3556 0 -1 305
box -2 -3 10 103
use FILL  FILL_3_2
timestamp 1696145522
transform -1 0 3564 0 -1 305
box -2 -3 10 103
use BUFX4  BUFX4_136
timestamp 1696145522
transform 1 0 4 0 1 305
box -2 -3 34 103
use BUFX4  BUFX4_129
timestamp 1696145522
transform 1 0 36 0 1 305
box -2 -3 34 103
use BUFX4  BUFX4_137
timestamp 1696145522
transform 1 0 68 0 1 305
box -2 -3 34 103
use BUFX4  BUFX4_36
timestamp 1696145522
transform 1 0 100 0 1 305
box -2 -3 34 103
use BUFX4  BUFX4_192
timestamp 1696145522
transform 1 0 132 0 1 305
box -2 -3 34 103
use BUFX4  BUFX4_195
timestamp 1696145522
transform 1 0 164 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_56
timestamp 1696145522
transform 1 0 196 0 1 305
box -2 -3 34 103
use BUFX4  BUFX4_117
timestamp 1696145522
transform 1 0 228 0 1 305
box -2 -3 34 103
use BUFX4  BUFX4_37
timestamp 1696145522
transform 1 0 260 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_165
timestamp 1696145522
transform 1 0 292 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_121
timestamp 1696145522
transform -1 0 348 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_253
timestamp 1696145522
transform -1 0 380 0 1 305
box -2 -3 34 103
use INVX1  INVX1_102
timestamp 1696145522
transform -1 0 396 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_279
timestamp 1696145522
transform -1 0 428 0 1 305
box -2 -3 34 103
use INVX1  INVX1_122
timestamp 1696145522
transform -1 0 444 0 1 305
box -2 -3 18 103
use MUX2X1  MUX2X1_2
timestamp 1696145522
transform -1 0 492 0 1 305
box -2 -3 50 103
use FILL  FILL_3_0_0
timestamp 1696145522
transform -1 0 500 0 1 305
box -2 -3 10 103
use FILL  FILL_3_0_1
timestamp 1696145522
transform -1 0 508 0 1 305
box -2 -3 10 103
use OAI21X1  OAI21X1_192
timestamp 1696145522
transform -1 0 540 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_563
timestamp 1696145522
transform 1 0 540 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_686
timestamp 1696145522
transform -1 0 596 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_298
timestamp 1696145522
transform 1 0 596 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_297
timestamp 1696145522
transform -1 0 660 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_687
timestamp 1696145522
transform -1 0 692 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_126
timestamp 1696145522
transform -1 0 716 0 1 305
box -2 -3 26 103
use INVX1  INVX1_288
timestamp 1696145522
transform -1 0 732 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_717
timestamp 1696145522
transform 1 0 732 0 1 305
box -2 -3 34 103
use MUX2X1  MUX2X1_110
timestamp 1696145522
transform 1 0 764 0 1 305
box -2 -3 50 103
use MUX2X1  MUX2X1_76
timestamp 1696145522
transform 1 0 812 0 1 305
box -2 -3 50 103
use NAND2X1  NAND2X1_580
timestamp 1696145522
transform -1 0 884 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_720
timestamp 1696145522
transform -1 0 916 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_721
timestamp 1696145522
transform -1 0 948 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_112
timestamp 1696145522
transform -1 0 980 0 1 305
box -2 -3 34 103
use INVX1  INVX1_101
timestamp 1696145522
transform -1 0 996 0 1 305
box -2 -3 18 103
use FILL  FILL_3_1_0
timestamp 1696145522
transform 1 0 996 0 1 305
box -2 -3 10 103
use FILL  FILL_3_1_1
timestamp 1696145522
transform 1 0 1004 0 1 305
box -2 -3 10 103
use MUX2X1  MUX2X1_88
timestamp 1696145522
transform 1 0 1012 0 1 305
box -2 -3 50 103
use MUX2X1  MUX2X1_90
timestamp 1696145522
transform 1 0 1060 0 1 305
box -2 -3 50 103
use MUX2X1  MUX2X1_100
timestamp 1696145522
transform 1 0 1108 0 1 305
box -2 -3 50 103
use MUX2X1  MUX2X1_98
timestamp 1696145522
transform 1 0 1156 0 1 305
box -2 -3 50 103
use MUX2X1  MUX2X1_93
timestamp 1696145522
transform 1 0 1204 0 1 305
box -2 -3 50 103
use NAND2X1  NAND2X1_163
timestamp 1696145522
transform -1 0 1276 0 1 305
box -2 -3 26 103
use MUX2X1  MUX2X1_86
timestamp 1696145522
transform 1 0 1276 0 1 305
box -2 -3 50 103
use MUX2X1  MUX2X1_97
timestamp 1696145522
transform 1 0 1324 0 1 305
box -2 -3 50 103
use OAI21X1  OAI21X1_110
timestamp 1696145522
transform -1 0 1404 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_70
timestamp 1696145522
transform 1 0 1404 0 1 305
box -2 -3 26 103
use INVX2  INVX2_11
timestamp 1696145522
transform -1 0 1444 0 1 305
box -2 -3 18 103
use NOR2X1  NOR2X1_55
timestamp 1696145522
transform -1 0 1468 0 1 305
box -2 -3 26 103
use INVX2  INVX2_10
timestamp 1696145522
transform 1 0 1468 0 1 305
box -2 -3 18 103
use BUFX4  BUFX4_178
timestamp 1696145522
transform 1 0 1484 0 1 305
box -2 -3 34 103
use FILL  FILL_3_2_0
timestamp 1696145522
transform -1 0 1524 0 1 305
box -2 -3 10 103
use FILL  FILL_3_2_1
timestamp 1696145522
transform -1 0 1532 0 1 305
box -2 -3 10 103
use INVX2  INVX2_14
timestamp 1696145522
transform -1 0 1548 0 1 305
box -2 -3 18 103
use XOR2X1  XOR2X1_7
timestamp 1696145522
transform 1 0 1548 0 1 305
box -2 -3 58 103
use NOR2X1  NOR2X1_17
timestamp 1696145522
transform -1 0 1628 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_741
timestamp 1696145522
transform 1 0 1628 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_730
timestamp 1696145522
transform -1 0 1692 0 1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_6
timestamp 1696145522
transform -1 0 1724 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_428
timestamp 1696145522
transform 1 0 1724 0 1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_308
timestamp 1696145522
transform 1 0 1748 0 1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_7
timestamp 1696145522
transform 1 0 1780 0 1 305
box -2 -3 34 103
use AOI22X1  AOI22X1_33
timestamp 1696145522
transform -1 0 1852 0 1 305
box -2 -3 42 103
use NOR2X1  NOR2X1_409
timestamp 1696145522
transform -1 0 1876 0 1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_24
timestamp 1696145522
transform 1 0 1876 0 1 305
box -2 -3 26 103
use NOR2X1  NOR2X1_22
timestamp 1696145522
transform -1 0 1924 0 1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_25
timestamp 1696145522
transform 1 0 1924 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_756
timestamp 1696145522
transform 1 0 1948 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_57
timestamp 1696145522
transform -1 0 2004 0 1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_196
timestamp 1696145522
transform -1 0 2028 0 1 305
box -2 -3 26 103
use FILL  FILL_3_3_0
timestamp 1696145522
transform -1 0 2036 0 1 305
box -2 -3 10 103
use FILL  FILL_3_3_1
timestamp 1696145522
transform -1 0 2044 0 1 305
box -2 -3 10 103
use OAI21X1  OAI21X1_750
timestamp 1696145522
transform -1 0 2076 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_195
timestamp 1696145522
transform -1 0 2100 0 1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_24
timestamp 1696145522
transform 1 0 2100 0 1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_61
timestamp 1696145522
transform -1 0 2164 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_23
timestamp 1696145522
transform 1 0 2164 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_11
timestamp 1696145522
transform 1 0 2188 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_751
timestamp 1696145522
transform 1 0 2220 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_24
timestamp 1696145522
transform -1 0 2276 0 1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_9
timestamp 1696145522
transform 1 0 2276 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_14
timestamp 1696145522
transform 1 0 2308 0 1 305
box -2 -3 34 103
use INVX1  INVX1_303
timestamp 1696145522
transform 1 0 2340 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_777
timestamp 1696145522
transform -1 0 2388 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_782
timestamp 1696145522
transform 1 0 2388 0 1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_326
timestamp 1696145522
transform 1 0 2420 0 1 305
box -2 -3 34 103
use INVX2  INVX2_22
timestamp 1696145522
transform -1 0 2468 0 1 305
box -2 -3 18 103
use INVX2  INVX2_16
timestamp 1696145522
transform 1 0 2468 0 1 305
box -2 -3 18 103
use INVX1  INVX1_305
timestamp 1696145522
transform 1 0 2484 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_794
timestamp 1696145522
transform 1 0 2500 0 1 305
box -2 -3 34 103
use FILL  FILL_3_4_0
timestamp 1696145522
transform 1 0 2532 0 1 305
box -2 -3 10 103
use FILL  FILL_3_4_1
timestamp 1696145522
transform 1 0 2540 0 1 305
box -2 -3 10 103
use AOI21X1  AOI21X1_10
timestamp 1696145522
transform 1 0 2548 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_153
timestamp 1696145522
transform 1 0 2580 0 1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_12
timestamp 1696145522
transform -1 0 2644 0 1 305
box -2 -3 34 103
use AOI22X1  AOI22X1_43
timestamp 1696145522
transform -1 0 2684 0 1 305
box -2 -3 42 103
use INVX1  INVX1_311
timestamp 1696145522
transform 1 0 2684 0 1 305
box -2 -3 18 103
use NAND3X1  NAND3X1_64
timestamp 1696145522
transform 1 0 2700 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_844
timestamp 1696145522
transform -1 0 2764 0 1 305
box -2 -3 34 103
use INVX1  INVX1_309
timestamp 1696145522
transform -1 0 2780 0 1 305
box -2 -3 18 103
use OAI21X1  OAI21X1_835
timestamp 1696145522
transform 1 0 2780 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_833
timestamp 1696145522
transform -1 0 2844 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_831
timestamp 1696145522
transform 1 0 2844 0 1 305
box -2 -3 34 103
use AOI21X1  AOI21X1_14
timestamp 1696145522
transform 1 0 2876 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_29
timestamp 1696145522
transform 1 0 2908 0 1 305
box -2 -3 26 103
use OAI21X1  OAI21X1_18
timestamp 1696145522
transform 1 0 2932 0 1 305
box -2 -3 34 103
use INVX1  INVX1_312
timestamp 1696145522
transform 1 0 2964 0 1 305
box -2 -3 18 103
use AOI21X1  AOI21X1_351
timestamp 1696145522
transform -1 0 3012 0 1 305
box -2 -3 34 103
use NAND3X1  NAND3X1_1
timestamp 1696145522
transform -1 0 3044 0 1 305
box -2 -3 34 103
use FILL  FILL_3_5_0
timestamp 1696145522
transform 1 0 3044 0 1 305
box -2 -3 10 103
use FILL  FILL_3_5_1
timestamp 1696145522
transform 1 0 3052 0 1 305
box -2 -3 10 103
use AOI22X1  AOI22X1_44
timestamp 1696145522
transform 1 0 3060 0 1 305
box -2 -3 42 103
use AOI21X1  AOI21X1_13
timestamp 1696145522
transform -1 0 3132 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_832
timestamp 1696145522
transform 1 0 3132 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_17
timestamp 1696145522
transform 1 0 3164 0 1 305
box -2 -3 34 103
use OAI21X1  OAI21X1_15
timestamp 1696145522
transform 1 0 3196 0 1 305
box -2 -3 34 103
use NAND2X1  NAND2X1_32
timestamp 1696145522
transform 1 0 3228 0 1 305
box -2 -3 26 103
use INVX2  INVX2_19
timestamp 1696145522
transform -1 0 3268 0 1 305
box -2 -3 18 103
use NAND2X1  NAND2X1_33
timestamp 1696145522
transform -1 0 3292 0 1 305
box -2 -3 26 103
use NOR2X1  NOR2X1_40
timestamp 1696145522
transform -1 0 3316 0 1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_31
timestamp 1696145522
transform -1 0 3340 0 1 305
box -2 -3 26 103
use INVX1  INVX1_16
timestamp 1696145522
transform -1 0 3356 0 1 305
box -2 -3 18 103
use NOR2X1  NOR2X1_476
timestamp 1696145522
transform 1 0 3356 0 1 305
box -2 -3 26 103
use AOI22X1  AOI22X1_41
timestamp 1696145522
transform 1 0 3380 0 1 305
box -2 -3 42 103
use AOI21X1  AOI21X1_352
timestamp 1696145522
transform -1 0 3452 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_472
timestamp 1696145522
transform -1 0 3476 0 1 305
box -2 -3 26 103
use INVX1  INVX1_313
timestamp 1696145522
transform 1 0 3476 0 1 305
box -2 -3 18 103
use NOR2X1  NOR2X1_35
timestamp 1696145522
transform 1 0 3492 0 1 305
box -2 -3 26 103
use AOI21X1  AOI21X1_11
timestamp 1696145522
transform 1 0 3516 0 1 305
box -2 -3 34 103
use FILL  FILL_4_1
timestamp 1696145522
transform 1 0 3548 0 1 305
box -2 -3 10 103
use FILL  FILL_4_2
timestamp 1696145522
transform 1 0 3556 0 1 305
box -2 -3 10 103
use INVX8  INVX8_3
timestamp 1696145522
transform -1 0 44 0 -1 505
box -2 -3 42 103
use BUFX4  BUFX4_133
timestamp 1696145522
transform 1 0 44 0 -1 505
box -2 -3 34 103
use INVX1  INVX1_36
timestamp 1696145522
transform -1 0 92 0 -1 505
box -2 -3 18 103
use BUFX4  BUFX4_135
timestamp 1696145522
transform 1 0 92 0 -1 505
box -2 -3 34 103
use BUFX4  BUFX4_34
timestamp 1696145522
transform 1 0 124 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_188
timestamp 1696145522
transform 1 0 156 0 -1 505
box -2 -3 34 103
use INVX1  INVX1_89
timestamp 1696145522
transform 1 0 188 0 -1 505
box -2 -3 18 103
use NAND2X1  NAND2X1_108
timestamp 1696145522
transform 1 0 204 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_189
timestamp 1696145522
transform 1 0 228 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_97
timestamp 1696145522
transform -1 0 292 0 -1 505
box -2 -3 34 103
use INVX1  INVX1_58
timestamp 1696145522
transform -1 0 308 0 -1 505
box -2 -3 18 103
use INVX1  INVX1_59
timestamp 1696145522
transform 1 0 308 0 -1 505
box -2 -3 18 103
use NAND2X1  NAND2X1_303
timestamp 1696145522
transform 1 0 324 0 -1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_240
timestamp 1696145522
transform 1 0 348 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_208
timestamp 1696145522
transform -1 0 404 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_239
timestamp 1696145522
transform 1 0 404 0 -1 505
box -2 -3 26 103
use BUFX4  BUFX4_123
timestamp 1696145522
transform 1 0 428 0 -1 505
box -2 -3 34 103
use BUFX4  BUFX4_125
timestamp 1696145522
transform 1 0 460 0 -1 505
box -2 -3 34 103
use FILL  FILL_4_0_0
timestamp 1696145522
transform 1 0 492 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_0_1
timestamp 1696145522
transform 1 0 500 0 -1 505
box -2 -3 10 103
use NAND2X1  NAND2X1_576
timestamp 1696145522
transform 1 0 508 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_716
timestamp 1696145522
transform -1 0 564 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_36
timestamp 1696145522
transform -1 0 596 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_86
timestamp 1696145522
transform -1 0 620 0 -1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_602
timestamp 1696145522
transform 1 0 620 0 -1 505
box -2 -3 26 103
use INVX1  INVX1_291
timestamp 1696145522
transform 1 0 644 0 -1 505
box -2 -3 18 103
use NAND2X1  NAND2X1_564
timestamp 1696145522
transform 1 0 660 0 -1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_595
timestamp 1696145522
transform 1 0 684 0 -1 505
box -2 -3 26 103
use INVX1  INVX1_287
timestamp 1696145522
transform 1 0 708 0 -1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_688
timestamp 1696145522
transform 1 0 724 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_578
timestamp 1696145522
transform 1 0 756 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_718
timestamp 1696145522
transform 1 0 780 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_159
timestamp 1696145522
transform -1 0 836 0 -1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_425
timestamp 1696145522
transform -1 0 860 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_212
timestamp 1696145522
transform -1 0 892 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_315
timestamp 1696145522
transform 1 0 892 0 -1 505
box -2 -3 34 103
use INVX1  INVX1_103
timestamp 1696145522
transform 1 0 924 0 -1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_314
timestamp 1696145522
transform -1 0 972 0 -1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_131
timestamp 1696145522
transform -1 0 996 0 -1 505
box -2 -3 26 103
use FILL  FILL_4_1_0
timestamp 1696145522
transform -1 0 1004 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_1_1
timestamp 1696145522
transform -1 0 1012 0 -1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_95
timestamp 1696145522
transform -1 0 1044 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_140
timestamp 1696145522
transform -1 0 1068 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_693
timestamp 1696145522
transform 1 0 1068 0 -1 505
box -2 -3 34 103
use MUX2X1  MUX2X1_81
timestamp 1696145522
transform 1 0 1100 0 -1 505
box -2 -3 50 103
use MUX2X1  MUX2X1_83
timestamp 1696145522
transform 1 0 1148 0 -1 505
box -2 -3 50 103
use MUX2X1  MUX2X1_94
timestamp 1696145522
transform 1 0 1196 0 -1 505
box -2 -3 50 103
use MUX2X1  MUX2X1_87
timestamp 1696145522
transform 1 0 1244 0 -1 505
box -2 -3 50 103
use MUX2X1  MUX2X1_108
timestamp 1696145522
transform 1 0 1292 0 -1 505
box -2 -3 50 103
use XOR2X1  XOR2X1_4
timestamp 1696145522
transform 1 0 1340 0 -1 505
box -2 -3 58 103
use OAI21X1  OAI21X1_701
timestamp 1696145522
transform 1 0 1396 0 -1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_16
timestamp 1696145522
transform 1 0 1428 0 -1 505
box -2 -3 26 103
use BUFX4  BUFX4_181
timestamp 1696145522
transform -1 0 1484 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_731
timestamp 1696145522
transform 1 0 1484 0 -1 505
box -2 -3 34 103
use FILL  FILL_4_2_0
timestamp 1696145522
transform 1 0 1516 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_2_1
timestamp 1696145522
transform 1 0 1524 0 -1 505
box -2 -3 10 103
use BUFX4  BUFX4_109
timestamp 1696145522
transform 1 0 1532 0 -1 505
box -2 -3 34 103
use INVX1  INVX1_289
timestamp 1696145522
transform 1 0 1564 0 -1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_702
timestamp 1696145522
transform -1 0 1612 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_742
timestamp 1696145522
transform 1 0 1612 0 -1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_311
timestamp 1696145522
transform 1 0 1644 0 -1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_301
timestamp 1696145522
transform -1 0 1708 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_700
timestamp 1696145522
transform 1 0 1708 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_567
timestamp 1696145522
transform 1 0 1740 0 -1 505
box -2 -3 26 103
use NAND3X1  NAND3X1_57
timestamp 1696145522
transform -1 0 1796 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_697
timestamp 1696145522
transform 1 0 1796 0 -1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_299
timestamp 1696145522
transform -1 0 1860 0 -1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_443
timestamp 1696145522
transform -1 0 1884 0 -1 505
box -2 -3 26 103
use INVX1  INVX1_301
timestamp 1696145522
transform 1 0 1884 0 -1 505
box -2 -3 18 103
use NAND3X1  NAND3X1_60
timestamp 1696145522
transform -1 0 1932 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_73
timestamp 1696145522
transform 1 0 1932 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_12
timestamp 1696145522
transform -1 0 1988 0 -1 505
box -2 -3 34 103
use AOI22X1  AOI22X1_35
timestamp 1696145522
transform -1 0 2028 0 -1 505
box -2 -3 42 103
use FILL  FILL_4_3_0
timestamp 1696145522
transform -1 0 2036 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_3_1
timestamp 1696145522
transform -1 0 2044 0 -1 505
box -2 -3 10 103
use INVX1  INVX1_297
timestamp 1696145522
transform -1 0 2060 0 -1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_778
timestamp 1696145522
transform -1 0 2092 0 -1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_439
timestamp 1696145522
transform -1 0 2116 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_775
timestamp 1696145522
transform -1 0 2148 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_13
timestamp 1696145522
transform -1 0 2180 0 -1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_321
timestamp 1696145522
transform 1 0 2180 0 -1 505
box -2 -3 34 103
use OR2X2  OR2X2_41
timestamp 1696145522
transform -1 0 2244 0 -1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_323
timestamp 1696145522
transform 1 0 2244 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_779
timestamp 1696145522
transform -1 0 2308 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_776
timestamp 1696145522
transform -1 0 2340 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_781
timestamp 1696145522
transform 1 0 2340 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_799
timestamp 1696145522
transform -1 0 2404 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_604
timestamp 1696145522
transform -1 0 2428 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_793
timestamp 1696145522
transform -1 0 2460 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_804
timestamp 1696145522
transform 1 0 2460 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_795
timestamp 1696145522
transform 1 0 2492 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_622
timestamp 1696145522
transform -1 0 2548 0 -1 505
box -2 -3 26 103
use FILL  FILL_4_4_0
timestamp 1696145522
transform -1 0 2556 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_4_1
timestamp 1696145522
transform -1 0 2564 0 -1 505
box -2 -3 10 103
use AOI21X1  AOI21X1_347
timestamp 1696145522
transform -1 0 2596 0 -1 505
box -2 -3 34 103
use INVX2  INVX2_17
timestamp 1696145522
transform 1 0 2596 0 -1 505
box -2 -3 18 103
use AOI21X1  AOI21X1_333
timestamp 1696145522
transform 1 0 2612 0 -1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_457
timestamp 1696145522
transform -1 0 2668 0 -1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_109
timestamp 1696145522
transform 1 0 2668 0 -1 505
box -2 -3 26 103
use NAND3X1  NAND3X1_65
timestamp 1696145522
transform 1 0 2692 0 -1 505
box -2 -3 34 103
use INVX1  INVX1_306
timestamp 1696145522
transform 1 0 2724 0 -1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_807
timestamp 1696145522
transform -1 0 2772 0 -1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_332
timestamp 1696145522
transform -1 0 2804 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_811
timestamp 1696145522
transform 1 0 2804 0 -1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_463
timestamp 1696145522
transform 1 0 2836 0 -1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_459
timestamp 1696145522
transform 1 0 2860 0 -1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_613
timestamp 1696145522
transform 1 0 2884 0 -1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_614
timestamp 1696145522
transform -1 0 2932 0 -1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_824
timestamp 1696145522
transform -1 0 2964 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_819
timestamp 1696145522
transform -1 0 2996 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_626
timestamp 1696145522
transform -1 0 3020 0 -1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_363
timestamp 1696145522
transform -1 0 3052 0 -1 505
box -2 -3 34 103
use FILL  FILL_4_5_0
timestamp 1696145522
transform 1 0 3052 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_5_1
timestamp 1696145522
transform 1 0 3060 0 -1 505
box -2 -3 10 103
use INVX2  INVX2_93
timestamp 1696145522
transform 1 0 3068 0 -1 505
box -2 -3 18 103
use AOI21X1  AOI21X1_337
timestamp 1696145522
transform 1 0 3084 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_851
timestamp 1696145522
transform -1 0 3148 0 -1 505
box -2 -3 34 103
use INVX2  INVX2_18
timestamp 1696145522
transform -1 0 3164 0 -1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_858
timestamp 1696145522
transform 1 0 3164 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_618
timestamp 1696145522
transform -1 0 3220 0 -1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_340
timestamp 1696145522
transform -1 0 3252 0 -1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_360
timestamp 1696145522
transform -1 0 3284 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_857
timestamp 1696145522
transform -1 0 3316 0 -1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_338
timestamp 1696145522
transform 1 0 3316 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_823
timestamp 1696145522
transform -1 0 3380 0 -1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_856
timestamp 1696145522
transform -1 0 3412 0 -1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_359
timestamp 1696145522
transform -1 0 3444 0 -1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_15
timestamp 1696145522
transform 1 0 3444 0 -1 505
box -2 -3 98 103
use INVX2  INVX2_94
timestamp 1696145522
transform 1 0 3540 0 -1 505
box -2 -3 18 103
use FILL  FILL_5_1
timestamp 1696145522
transform -1 0 3564 0 -1 505
box -2 -3 10 103
use BUFX4  BUFX4_128
timestamp 1696145522
transform 1 0 4 0 1 505
box -2 -3 34 103
use BUFX4  BUFX4_132
timestamp 1696145522
transform 1 0 36 0 1 505
box -2 -3 34 103
use BUFX4  BUFX4_134
timestamp 1696145522
transform 1 0 68 0 1 505
box -2 -3 34 103
use BUFX4  BUFX4_33
timestamp 1696145522
transform 1 0 100 0 1 505
box -2 -3 34 103
use BUFX4  BUFX4_40
timestamp 1696145522
transform 1 0 132 0 1 505
box -2 -3 34 103
use BUFX4  BUFX4_39
timestamp 1696145522
transform 1 0 164 0 1 505
box -2 -3 34 103
use INVX1  INVX1_45
timestamp 1696145522
transform -1 0 212 0 1 505
box -2 -3 18 103
use BUFX4  BUFX4_131
timestamp 1696145522
transform 1 0 212 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_247
timestamp 1696145522
transform 1 0 244 0 1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_142
timestamp 1696145522
transform -1 0 292 0 1 505
box -2 -3 26 103
use BUFX4  BUFX4_38
timestamp 1696145522
transform 1 0 292 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_280
timestamp 1696145522
transform 1 0 324 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_209
timestamp 1696145522
transform 1 0 356 0 1 505
box -2 -3 34 103
use INVX1  INVX1_136
timestamp 1696145522
transform 1 0 388 0 1 505
box -2 -3 18 103
use INVX1  INVX1_123
timestamp 1696145522
transform 1 0 404 0 1 505
box -2 -3 18 103
use NAND2X1  NAND2X1_333
timestamp 1696145522
transform 1 0 420 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_444
timestamp 1696145522
transform 1 0 444 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_418
timestamp 1696145522
transform 1 0 476 0 1 505
box -2 -3 26 103
use FILL  FILL_5_0_0
timestamp 1696145522
transform 1 0 500 0 1 505
box -2 -3 10 103
use FILL  FILL_5_0_1
timestamp 1696145522
transform 1 0 508 0 1 505
box -2 -3 10 103
use NAND2X1  NAND2X1_559
timestamp 1696145522
transform 1 0 516 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_681
timestamp 1696145522
transform -1 0 572 0 1 505
box -2 -3 34 103
use INVX1  INVX1_285
timestamp 1696145522
transform -1 0 588 0 1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_679
timestamp 1696145522
transform -1 0 620 0 1 505
box -2 -3 34 103
use OR2X2  OR2X2_22
timestamp 1696145522
transform -1 0 652 0 1 505
box -2 -3 34 103
use MUX2X1  MUX2X1_106
timestamp 1696145522
transform 1 0 652 0 1 505
box -2 -3 50 103
use INVX1  INVX1_98
timestamp 1696145522
transform 1 0 700 0 1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_747
timestamp 1696145522
transform -1 0 748 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_603
timestamp 1696145522
transform 1 0 748 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_769
timestamp 1696145522
transform -1 0 804 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_418
timestamp 1696145522
transform 1 0 804 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_417
timestamp 1696145522
transform -1 0 868 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_115
timestamp 1696145522
transform 1 0 868 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_598
timestamp 1696145522
transform 1 0 900 0 1 505
box -2 -3 26 103
use MUX2X1  MUX2X1_96
timestamp 1696145522
transform 1 0 924 0 1 505
box -2 -3 50 103
use NOR2X1  NOR2X1_147
timestamp 1696145522
transform -1 0 996 0 1 505
box -2 -3 26 103
use FILL  FILL_5_1_0
timestamp 1696145522
transform 1 0 996 0 1 505
box -2 -3 10 103
use FILL  FILL_5_1_1
timestamp 1696145522
transform 1 0 1004 0 1 505
box -2 -3 10 103
use NAND2X1  NAND2X1_244
timestamp 1696145522
transform 1 0 1012 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_739
timestamp 1696145522
transform 1 0 1036 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_760
timestamp 1696145522
transform -1 0 1100 0 1 505
box -2 -3 34 103
use MUX2X1  MUX2X1_101
timestamp 1696145522
transform -1 0 1148 0 1 505
box -2 -3 50 103
use MUX2X1  MUX2X1_113
timestamp 1696145522
transform -1 0 1196 0 1 505
box -2 -3 50 103
use OAI21X1  OAI21X1_388
timestamp 1696145522
transform 1 0 1196 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_387
timestamp 1696145522
transform -1 0 1260 0 1 505
box -2 -3 34 103
use INVX1  INVX1_166
timestamp 1696145522
transform -1 0 1276 0 1 505
box -2 -3 18 103
use MUX2X1  MUX2X1_99
timestamp 1696145522
transform -1 0 1324 0 1 505
box -2 -3 50 103
use NAND3X1  NAND3X1_7
timestamp 1696145522
transform -1 0 1356 0 1 505
box -2 -3 34 103
use MUX2X1  MUX2X1_102
timestamp 1696145522
transform 1 0 1356 0 1 505
box -2 -3 50 103
use MUX2X1  MUX2X1_95
timestamp 1696145522
transform 1 0 1404 0 1 505
box -2 -3 50 103
use MUX2X1  MUX2X1_109
timestamp 1696145522
transform 1 0 1452 0 1 505
box -2 -3 50 103
use FILL  FILL_5_2_0
timestamp 1696145522
transform 1 0 1500 0 1 505
box -2 -3 10 103
use FILL  FILL_5_2_1
timestamp 1696145522
transform 1 0 1508 0 1 505
box -2 -3 10 103
use MUX2X1  MUX2X1_119
timestamp 1696145522
transform 1 0 1516 0 1 505
box -2 -3 50 103
use BUFX4  BUFX4_179
timestamp 1696145522
transform -1 0 1596 0 1 505
box -2 -3 34 103
use BUFX4  BUFX4_111
timestamp 1696145522
transform 1 0 1596 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_59
timestamp 1696145522
transform 1 0 1628 0 1 505
box -2 -3 34 103
use BUFX4  BUFX4_183
timestamp 1696145522
transform 1 0 1660 0 1 505
box -2 -3 34 103
use BUFX4  BUFX4_114
timestamp 1696145522
transform 1 0 1692 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_746
timestamp 1696145522
transform 1 0 1724 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_437
timestamp 1696145522
transform -1 0 1780 0 1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_594
timestamp 1696145522
transform -1 0 1804 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_745
timestamp 1696145522
transform -1 0 1836 0 1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_313
timestamp 1696145522
transform 1 0 1836 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_58
timestamp 1696145522
transform 1 0 1868 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_753
timestamp 1696145522
transform 1 0 1900 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_27
timestamp 1696145522
transform 1 0 1932 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_755
timestamp 1696145522
transform 1 0 1956 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_754
timestamp 1696145522
transform -1 0 2020 0 1 505
box -2 -3 34 103
use FILL  FILL_5_3_0
timestamp 1696145522
transform -1 0 2028 0 1 505
box -2 -3 10 103
use FILL  FILL_5_3_1
timestamp 1696145522
transform -1 0 2036 0 1 505
box -2 -3 10 103
use NOR2X1  NOR2X1_440
timestamp 1696145522
transform -1 0 2060 0 1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_597
timestamp 1696145522
transform 1 0 2060 0 1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_441
timestamp 1696145522
transform -1 0 2108 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_766
timestamp 1696145522
transform -1 0 2140 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_767
timestamp 1696145522
transform -1 0 2172 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_6
timestamp 1696145522
transform 1 0 2172 0 1 505
box -2 -3 98 103
use INVX1  INVX1_266
timestamp 1696145522
transform 1 0 2268 0 1 505
box -2 -3 18 103
use AOI22X1  AOI22X1_34
timestamp 1696145522
transform 1 0 2284 0 1 505
box -2 -3 42 103
use BUFX2  BUFX2_5
timestamp 1696145522
transform 1 0 2324 0 1 505
box -2 -3 26 103
use NAND3X1  NAND3X1_46
timestamp 1696145522
transform 1 0 2348 0 1 505
box -2 -3 34 103
use INVX1  INVX1_267
timestamp 1696145522
transform -1 0 2396 0 1 505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_5
timestamp 1696145522
transform -1 0 2492 0 1 505
box -2 -3 98 103
use AOI21X1  AOI21X1_327
timestamp 1696145522
transform -1 0 2524 0 1 505
box -2 -3 34 103
use FILL  FILL_5_4_0
timestamp 1696145522
transform 1 0 2524 0 1 505
box -2 -3 10 103
use FILL  FILL_5_4_1
timestamp 1696145522
transform 1 0 2532 0 1 505
box -2 -3 10 103
use OR2X2  OR2X2_42
timestamp 1696145522
transform 1 0 2540 0 1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_331
timestamp 1696145522
transform -1 0 2604 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_805
timestamp 1696145522
transform -1 0 2636 0 1 505
box -2 -3 34 103
use NAND3X1  NAND3X1_63
timestamp 1696145522
transform 1 0 2636 0 1 505
box -2 -3 34 103
use AOI22X1  AOI22X1_37
timestamp 1696145522
transform 1 0 2668 0 1 505
box -2 -3 42 103
use INVX1  INVX1_17
timestamp 1696145522
transform 1 0 2708 0 1 505
box -2 -3 18 103
use NAND3X1  NAND3X1_2
timestamp 1696145522
transform 1 0 2724 0 1 505
box -2 -3 34 103
use BUFX2  BUFX2_10
timestamp 1696145522
transform 1 0 2756 0 1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_454
timestamp 1696145522
transform 1 0 2780 0 1 505
box -2 -3 26 103
use OR2X2  OR2X2_1
timestamp 1696145522
transform 1 0 2804 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_19
timestamp 1696145522
transform 1 0 2836 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_822
timestamp 1696145522
transform 1 0 2868 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_460
timestamp 1696145522
transform 1 0 2900 0 1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_28
timestamp 1696145522
transform -1 0 2948 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_820
timestamp 1696145522
transform 1 0 2948 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_855
timestamp 1696145522
transform 1 0 2980 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_624
timestamp 1696145522
transform -1 0 3036 0 1 505
box -2 -3 26 103
use FILL  FILL_5_5_0
timestamp 1696145522
transform -1 0 3044 0 1 505
box -2 -3 10 103
use FILL  FILL_5_5_1
timestamp 1696145522
transform -1 0 3052 0 1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_854
timestamp 1696145522
transform -1 0 3084 0 1 505
box -2 -3 34 103
use INVX1  INVX1_307
timestamp 1696145522
transform -1 0 3100 0 1 505
box -2 -3 18 103
use NAND3X1  NAND3X1_67
timestamp 1696145522
transform 1 0 3100 0 1 505
box -2 -3 34 103
use OR2X2  OR2X2_45
timestamp 1696145522
transform -1 0 3164 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_479
timestamp 1696145522
transform -1 0 3188 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_361
timestamp 1696145522
transform 1 0 3188 0 1 505
box -2 -3 34 103
use OAI21X1  OAI21X1_859
timestamp 1696145522
transform 1 0 3220 0 1 505
box -2 -3 34 103
use INVX8  INVX8_19
timestamp 1696145522
transform -1 0 3292 0 1 505
box -2 -3 42 103
use AOI21X1  AOI21X1_365
timestamp 1696145522
transform 1 0 3292 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_480
timestamp 1696145522
transform 1 0 3324 0 1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_402
timestamp 1696145522
transform 1 0 3348 0 1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_625
timestamp 1696145522
transform 1 0 3372 0 1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_16
timestamp 1696145522
transform 1 0 3396 0 1 505
box -2 -3 98 103
use BUFX2  BUFX2_18
timestamp 1696145522
transform 1 0 3492 0 1 505
box -2 -3 26 103
use BUFX2  BUFX2_17
timestamp 1696145522
transform 1 0 3516 0 1 505
box -2 -3 26 103
use INVX2  INVX2_28
timestamp 1696145522
transform 1 0 3540 0 1 505
box -2 -3 18 103
use FILL  FILL_6_1
timestamp 1696145522
transform 1 0 3556 0 1 505
box -2 -3 10 103
use BUFX4  BUFX4_119
timestamp 1696145522
transform -1 0 36 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_87
timestamp 1696145522
transform 1 0 36 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_38
timestamp 1696145522
transform -1 0 92 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_278
timestamp 1696145522
transform 1 0 92 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_254
timestamp 1696145522
transform -1 0 148 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_309
timestamp 1696145522
transform 1 0 148 0 -1 705
box -2 -3 26 103
use BUFX4  BUFX4_42
timestamp 1696145522
transform 1 0 172 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_59
timestamp 1696145522
transform 1 0 204 0 -1 705
box -2 -3 34 103
use BUFX4  BUFX4_41
timestamp 1696145522
transform 1 0 236 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_215
timestamp 1696145522
transform -1 0 300 0 -1 705
box -2 -3 34 103
use BUFX4  BUFX4_127
timestamp 1696145522
transform 1 0 300 0 -1 705
box -2 -3 34 103
use BUFX4  BUFX4_20
timestamp 1696145522
transform 1 0 332 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_332
timestamp 1696145522
transform 1 0 364 0 -1 705
box -2 -3 26 103
use INVX1  INVX1_149
timestamp 1696145522
transform 1 0 388 0 -1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_319
timestamp 1696145522
transform 1 0 404 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_248
timestamp 1696145522
transform 1 0 436 0 -1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_166
timestamp 1696145522
transform -1 0 484 0 -1 705
box -2 -3 26 103
use FILL  FILL_6_0_0
timestamp 1696145522
transform -1 0 492 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_0_1
timestamp 1696145522
transform -1 0 500 0 -1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_320
timestamp 1696145522
transform -1 0 532 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_60
timestamp 1696145522
transform -1 0 564 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_380
timestamp 1696145522
transform 1 0 564 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_37
timestamp 1696145522
transform -1 0 620 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_429
timestamp 1696145522
transform -1 0 652 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_226
timestamp 1696145522
transform -1 0 676 0 -1 705
box -2 -3 26 103
use BUFX4  BUFX4_26
timestamp 1696145522
transform 1 0 676 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_159
timestamp 1696145522
transform -1 0 732 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_768
timestamp 1696145522
transform -1 0 764 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_573
timestamp 1696145522
transform 1 0 764 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_711
timestamp 1696145522
transform -1 0 820 0 -1 705
box -2 -3 34 103
use INVX1  INVX1_290
timestamp 1696145522
transform -1 0 836 0 -1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_369
timestamp 1696145522
transform 1 0 836 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_368
timestamp 1696145522
transform -1 0 900 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_127
timestamp 1696145522
transform -1 0 924 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_710
timestamp 1696145522
transform -1 0 956 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_814
timestamp 1696145522
transform -1 0 988 0 -1 705
box -2 -3 34 103
use FILL  FILL_6_1_0
timestamp 1696145522
transform 1 0 988 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_1_1
timestamp 1696145522
transform 1 0 996 0 -1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_213
timestamp 1696145522
transform 1 0 1004 0 -1 705
box -2 -3 34 103
use INVX1  INVX1_99
timestamp 1696145522
transform 1 0 1036 0 -1 705
box -2 -3 18 103
use NAND2X1  NAND2X1_593
timestamp 1696145522
transform -1 0 1076 0 -1 705
box -2 -3 26 103
use OR2X2  OR2X2_39
timestamp 1696145522
transform 1 0 1076 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_737
timestamp 1696145522
transform -1 0 1140 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_541
timestamp 1696145522
transform 1 0 1140 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_540
timestamp 1696145522
transform -1 0 1204 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_709
timestamp 1696145522
transform 1 0 1204 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_565
timestamp 1696145522
transform -1 0 1260 0 -1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_470
timestamp 1696145522
transform 1 0 1260 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_738
timestamp 1696145522
transform -1 0 1316 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_616
timestamp 1696145522
transform -1 0 1340 0 -1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_166
timestamp 1696145522
transform -1 0 1364 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_827
timestamp 1696145522
transform -1 0 1396 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_96
timestamp 1696145522
transform -1 0 1428 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_740
timestamp 1696145522
transform 1 0 1428 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_310
timestamp 1696145522
transform -1 0 1492 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_575
timestamp 1696145522
transform 1 0 1492 0 -1 705
box -2 -3 26 103
use FILL  FILL_6_2_0
timestamp 1696145522
transform -1 0 1524 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_2_1
timestamp 1696145522
transform -1 0 1532 0 -1 705
box -2 -3 10 103
use NOR2X1  NOR2X1_455
timestamp 1696145522
transform -1 0 1556 0 -1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_456
timestamp 1696145522
transform -1 0 1580 0 -1 705
box -2 -3 26 103
use BUFX4  BUFX4_180
timestamp 1696145522
transform -1 0 1612 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_438
timestamp 1696145522
transform 1 0 1612 0 -1 705
box -2 -3 26 103
use BUFX4  BUFX4_182
timestamp 1696145522
transform 1 0 1636 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_712
timestamp 1696145522
transform 1 0 1668 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_305
timestamp 1696145522
transform 1 0 1700 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_714
timestamp 1696145522
transform -1 0 1764 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_303
timestamp 1696145522
transform -1 0 1796 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_369
timestamp 1696145522
transform 1 0 1796 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_474
timestamp 1696145522
transform -1 0 1852 0 -1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_433
timestamp 1696145522
transform -1 0 1876 0 -1 705
box -2 -3 26 103
use BUFX4  BUFX4_113
timestamp 1696145522
transform 1 0 1876 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_451
timestamp 1696145522
transform 1 0 1908 0 -1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_330
timestamp 1696145522
transform -1 0 1956 0 -1 705
box -2 -3 26 103
use XNOR2X1  XNOR2X1_21
timestamp 1696145522
transform -1 0 2012 0 -1 705
box -2 -3 58 103
use NAND2X1  NAND2X1_608
timestamp 1696145522
transform -1 0 2036 0 -1 705
box -2 -3 26 103
use FILL  FILL_6_3_0
timestamp 1696145522
transform -1 0 2044 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_3_1
timestamp 1696145522
transform -1 0 2052 0 -1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_696
timestamp 1696145522
transform -1 0 2084 0 -1 705
box -2 -3 34 103
use AND2X2  AND2X2_51
timestamp 1696145522
transform 1 0 2084 0 -1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_62
timestamp 1696145522
transform -1 0 2148 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_429
timestamp 1696145522
transform -1 0 2172 0 -1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_314
timestamp 1696145522
transform 1 0 2172 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_434
timestamp 1696145522
transform 1 0 2204 0 -1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_4
timestamp 1696145522
transform 1 0 2228 0 -1 705
box -2 -3 98 103
use NOR2X1  NOR2X1_430
timestamp 1696145522
transform -1 0 2348 0 -1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_398
timestamp 1696145522
transform 1 0 2348 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_791
timestamp 1696145522
transform 1 0 2372 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_356
timestamp 1696145522
transform 1 0 2404 0 -1 705
box -2 -3 34 103
use AND2X2  AND2X2_65
timestamp 1696145522
transform 1 0 2436 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_792
timestamp 1696145522
transform -1 0 2500 0 -1 705
box -2 -3 34 103
use INVX1  INVX1_304
timestamp 1696145522
transform -1 0 2516 0 -1 705
box -2 -3 18 103
use FILL  FILL_6_4_0
timestamp 1696145522
transform 1 0 2516 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_4_1
timestamp 1696145522
transform 1 0 2524 0 -1 705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_8
timestamp 1696145522
transform 1 0 2532 0 -1 705
box -2 -3 98 103
use NOR2X1  NOR2X1_400
timestamp 1696145522
transform 1 0 2628 0 -1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_349
timestamp 1696145522
transform -1 0 2684 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_350
timestamp 1696145522
transform 1 0 2684 0 -1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_14
timestamp 1696145522
transform 1 0 2716 0 -1 705
box -2 -3 98 103
use AND2X2  AND2X2_58
timestamp 1696145522
transform 1 0 2812 0 -1 705
box -2 -3 34 103
use INVX2  INVX2_6
timestamp 1696145522
transform -1 0 2860 0 -1 705
box -2 -3 18 103
use BUFX4  BUFX4_14
timestamp 1696145522
transform -1 0 2892 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_821
timestamp 1696145522
transform 1 0 2892 0 -1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_339
timestamp 1696145522
transform -1 0 2956 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_825
timestamp 1696145522
transform -1 0 2988 0 -1 705
box -2 -3 34 103
use AOI22X1  AOI22X1_39
timestamp 1696145522
transform -1 0 3028 0 -1 705
box -2 -3 42 103
use NAND3X1  NAND3X1_68
timestamp 1696145522
transform -1 0 3060 0 -1 705
box -2 -3 34 103
use FILL  FILL_6_5_0
timestamp 1696145522
transform 1 0 3060 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_5_1
timestamp 1696145522
transform 1 0 3068 0 -1 705
box -2 -3 10 103
use AOI21X1  AOI21X1_334
timestamp 1696145522
transform 1 0 3076 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_812
timestamp 1696145522
transform 1 0 3108 0 -1 705
box -2 -3 34 103
use INVX1  INVX1_264
timestamp 1696145522
transform -1 0 3156 0 -1 705
box -2 -3 18 103
use AOI22X1  AOI22X1_40
timestamp 1696145522
transform -1 0 3196 0 -1 705
box -2 -3 42 103
use NAND3X1  NAND3X1_44
timestamp 1696145522
transform -1 0 3228 0 -1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_10
timestamp 1696145522
transform 1 0 3228 0 -1 705
box -2 -3 98 103
use INVX1  INVX1_263
timestamp 1696145522
transform -1 0 3340 0 -1 705
box -2 -3 18 103
use AOI22X1  AOI22X1_42
timestamp 1696145522
transform -1 0 3380 0 -1 705
box -2 -3 42 103
use BUFX4  BUFX4_11
timestamp 1696145522
transform -1 0 3412 0 -1 705
box -2 -3 34 103
use INVX1  INVX1_262
timestamp 1696145522
transform -1 0 3428 0 -1 705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_12
timestamp 1696145522
transform 1 0 3428 0 -1 705
box -2 -3 98 103
use BUFX2  BUFX2_12
timestamp 1696145522
transform 1 0 3524 0 -1 705
box -2 -3 26 103
use FILL  FILL_7_1
timestamp 1696145522
transform -1 0 3556 0 -1 705
box -2 -3 10 103
use FILL  FILL_7_2
timestamp 1696145522
transform -1 0 3564 0 -1 705
box -2 -3 10 103
use BUFX4  BUFX4_67
timestamp 1696145522
transform -1 0 36 0 1 705
box -2 -3 34 103
use INVX1  INVX1_91
timestamp 1696145522
transform 1 0 36 0 1 705
box -2 -3 18 103
use INVX1  INVX1_92
timestamp 1696145522
transform -1 0 68 0 1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_194
timestamp 1696145522
transform 1 0 68 0 1 705
box -2 -3 34 103
use INVX8  INVX8_2
timestamp 1696145522
transform -1 0 140 0 1 705
box -2 -3 42 103
use INVX1  INVX1_112
timestamp 1696145522
transform 1 0 140 0 1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_291
timestamp 1696145522
transform -1 0 188 0 1 705
box -2 -3 34 103
use INVX1  INVX1_37
timestamp 1696145522
transform 1 0 188 0 1 705
box -2 -3 18 103
use NAND2X1  NAND2X1_297
timestamp 1696145522
transform 1 0 204 0 1 705
box -2 -3 26 103
use INVX1  INVX1_46
timestamp 1696145522
transform 1 0 228 0 1 705
box -2 -3 18 103
use NAND2X1  NAND2X1_146
timestamp 1696145522
transform 1 0 244 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_100
timestamp 1696145522
transform -1 0 300 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_101
timestamp 1696145522
transform -1 0 332 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_145
timestamp 1696145522
transform 1 0 332 0 1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_361
timestamp 1696145522
transform 1 0 356 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_352
timestamp 1696145522
transform -1 0 412 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_281
timestamp 1696145522
transform 1 0 412 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_304
timestamp 1696145522
transform -1 0 468 0 1 705
box -2 -3 26 103
use INVX1  INVX1_137
timestamp 1696145522
transform 1 0 468 0 1 705
box -2 -3 18 103
use FILL  FILL_7_0_0
timestamp 1696145522
transform -1 0 492 0 1 705
box -2 -3 10 103
use FILL  FILL_7_0_1
timestamp 1696145522
transform -1 0 500 0 1 705
box -2 -3 10 103
use NAND2X1  NAND2X1_109
timestamp 1696145522
transform -1 0 524 0 1 705
box -2 -3 26 103
use MUX2X1  MUX2X1_31
timestamp 1696145522
transform -1 0 572 0 1 705
box -2 -3 50 103
use NAND2X1  NAND2X1_347
timestamp 1696145522
transform 1 0 572 0 1 705
box -2 -3 26 103
use INVX1  INVX1_138
timestamp 1696145522
transform -1 0 612 0 1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_680
timestamp 1696145522
transform 1 0 612 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_582
timestamp 1696145522
transform -1 0 668 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_723
timestamp 1696145522
transform -1 0 700 0 1 705
box -2 -3 34 103
use INVX1  INVX1_292
timestamp 1696145522
transform 1 0 700 0 1 705
box -2 -3 18 103
use INVX1  INVX1_177
timestamp 1696145522
transform 1 0 716 0 1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_397
timestamp 1696145522
transform 1 0 732 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_396
timestamp 1696145522
transform -1 0 796 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_583
timestamp 1696145522
transform 1 0 796 0 1 705
box -2 -3 26 103
use MUX2X1  MUX2X1_74
timestamp 1696145522
transform 1 0 820 0 1 705
box -2 -3 50 103
use NAND2X1  NAND2X1_591
timestamp 1696145522
transform 1 0 868 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_736
timestamp 1696145522
transform 1 0 892 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_574
timestamp 1696145522
transform -1 0 948 0 1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_612
timestamp 1696145522
transform -1 0 972 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_708
timestamp 1696145522
transform 1 0 972 0 1 705
box -2 -3 34 103
use FILL  FILL_7_1_0
timestamp 1696145522
transform -1 0 1012 0 1 705
box -2 -3 10 103
use FILL  FILL_7_1_1
timestamp 1696145522
transform -1 0 1020 0 1 705
box -2 -3 10 103
use NAND2X1  NAND2X1_600
timestamp 1696145522
transform -1 0 1044 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_762
timestamp 1696145522
transform -1 0 1076 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_601
timestamp 1696145522
transform -1 0 1100 0 1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_592
timestamp 1696145522
transform 1 0 1100 0 1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_471
timestamp 1696145522
transform -1 0 1148 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_122
timestamp 1696145522
transform -1 0 1180 0 1 705
box -2 -3 34 103
use INVX1  INVX1_66
timestamp 1696145522
transform 1 0 1180 0 1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_554
timestamp 1696145522
transform 1 0 1196 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_770
timestamp 1696145522
transform -1 0 1260 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_846
timestamp 1696145522
transform 1 0 1260 0 1 705
box -2 -3 34 103
use MUX2X1  MUX2X1_114
timestamp 1696145522
transform 1 0 1292 0 1 705
box -2 -3 50 103
use MUX2X1  MUX2X1_115
timestamp 1696145522
transform 1 0 1340 0 1 705
box -2 -3 50 103
use NAND3X1  NAND3X1_56
timestamp 1696145522
transform -1 0 1420 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_141
timestamp 1696145522
transform -1 0 1444 0 1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_285
timestamp 1696145522
transform -1 0 1468 0 1 705
box -2 -3 26 103
use NAND3X1  NAND3X1_14
timestamp 1696145522
transform -1 0 1500 0 1 705
box -2 -3 34 103
use INVX1  INVX1_132
timestamp 1696145522
transform 1 0 1500 0 1 705
box -2 -3 18 103
use FILL  FILL_7_2_0
timestamp 1696145522
transform 1 0 1516 0 1 705
box -2 -3 10 103
use FILL  FILL_7_2_1
timestamp 1696145522
transform 1 0 1524 0 1 705
box -2 -3 10 103
use INVX1  INVX1_318
timestamp 1696145522
transform 1 0 1532 0 1 705
box -2 -3 18 103
use BUFX4  BUFX4_185
timestamp 1696145522
transform 1 0 1548 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_828
timestamp 1696145522
transform 1 0 1580 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_141
timestamp 1696145522
transform 1 0 1612 0 1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_571
timestamp 1696145522
transform -1 0 1660 0 1 705
box -2 -3 26 103
use OR2X2  OR2X2_43
timestamp 1696145522
transform 1 0 1660 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_442
timestamp 1696145522
transform -1 0 1716 0 1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_319
timestamp 1696145522
transform -1 0 1748 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_436
timestamp 1696145522
transform 1 0 1748 0 1 705
box -2 -3 26 103
use BUFX4  BUFX4_184
timestamp 1696145522
transform 1 0 1772 0 1 705
box -2 -3 34 103
use INVX4  INVX4_6
timestamp 1696145522
transform -1 0 1828 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_801
timestamp 1696145522
transform 1 0 1828 0 1 705
box -2 -3 34 103
use BUFX4  BUFX4_112
timestamp 1696145522
transform 1 0 1860 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_607
timestamp 1696145522
transform 1 0 1892 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_790
timestamp 1696145522
transform -1 0 1948 0 1 705
box -2 -3 34 103
use OR2X2  OR2X2_40
timestamp 1696145522
transform 1 0 1948 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_765
timestamp 1696145522
transform 1 0 1980 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_606
timestamp 1696145522
transform -1 0 2036 0 1 705
box -2 -3 26 103
use FILL  FILL_7_3_0
timestamp 1696145522
transform 1 0 2036 0 1 705
box -2 -3 10 103
use FILL  FILL_7_3_1
timestamp 1696145522
transform 1 0 2044 0 1 705
box -2 -3 10 103
use INVX1  INVX1_300
timestamp 1696145522
transform 1 0 2052 0 1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_780
timestamp 1696145522
transform 1 0 2068 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_771
timestamp 1696145522
transform -1 0 2132 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_764
timestamp 1696145522
transform 1 0 2132 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_320
timestamp 1696145522
transform 1 0 2164 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_444
timestamp 1696145522
transform -1 0 2220 0 1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_324
timestamp 1696145522
transform 1 0 2220 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_322
timestamp 1696145522
transform 1 0 2252 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_309
timestamp 1696145522
transform 1 0 2284 0 1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_3
timestamp 1696145522
transform 1 0 2316 0 1 705
box -2 -3 98 103
use NOR2X1  NOR2X1_453
timestamp 1696145522
transform -1 0 2436 0 1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_610
timestamp 1696145522
transform 1 0 2436 0 1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_325
timestamp 1696145522
transform 1 0 2460 0 1 705
box -2 -3 34 103
use FILL  FILL_7_4_0
timestamp 1696145522
transform 1 0 2492 0 1 705
box -2 -3 10 103
use FILL  FILL_7_4_1
timestamp 1696145522
transform 1 0 2500 0 1 705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_7
timestamp 1696145522
transform 1 0 2508 0 1 705
box -2 -3 98 103
use NOR2X1  NOR2X1_445
timestamp 1696145522
transform -1 0 2628 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_802
timestamp 1696145522
transform 1 0 2628 0 1 705
box -2 -3 34 103
use XNOR2X1  XNOR2X1_24
timestamp 1696145522
transform -1 0 2716 0 1 705
box -2 -3 58 103
use NOR2X1  NOR2X1_469
timestamp 1696145522
transform 1 0 2716 0 1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_336
timestamp 1696145522
transform 1 0 2740 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_396
timestamp 1696145522
transform 1 0 2772 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_842
timestamp 1696145522
transform 1 0 2796 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_843
timestamp 1696145522
transform -1 0 2860 0 1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_13
timestamp 1696145522
transform 1 0 2860 0 1 705
box -2 -3 98 103
use INVX1  INVX1_308
timestamp 1696145522
transform -1 0 2972 0 1 705
box -2 -3 18 103
use AND2X2  AND2X2_60
timestamp 1696145522
transform 1 0 2972 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_358
timestamp 1696145522
transform -1 0 3036 0 1 705
box -2 -3 34 103
use FILL  FILL_7_5_0
timestamp 1696145522
transform 1 0 3036 0 1 705
box -2 -3 10 103
use FILL  FILL_7_5_1
timestamp 1696145522
transform 1 0 3044 0 1 705
box -2 -3 10 103
use OAI21X1  OAI21X1_864
timestamp 1696145522
transform 1 0 3052 0 1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_45
timestamp 1696145522
transform -1 0 3116 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_535
timestamp 1696145522
transform -1 0 3140 0 1 705
box -2 -3 26 103
use NOR2X1  NOR2X1_397
timestamp 1696145522
transform -1 0 3164 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_803
timestamp 1696145522
transform -1 0 3196 0 1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_395
timestamp 1696145522
transform 1 0 3196 0 1 705
box -2 -3 26 103
use INVX1  INVX1_265
timestamp 1696145522
transform -1 0 3236 0 1 705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_9
timestamp 1696145522
transform 1 0 3236 0 1 705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_11
timestamp 1696145522
transform 1 0 3332 0 1 705
box -2 -3 98 103
use BUFX2  BUFX2_11
timestamp 1696145522
transform 1 0 3428 0 1 705
box -2 -3 26 103
use BUFX2  BUFX2_16
timestamp 1696145522
transform 1 0 3452 0 1 705
box -2 -3 26 103
use BUFX2  BUFX2_15
timestamp 1696145522
transform 1 0 3476 0 1 705
box -2 -3 26 103
use BUFX2  BUFX2_9
timestamp 1696145522
transform 1 0 3500 0 1 705
box -2 -3 26 103
use BUFX2  BUFX2_14
timestamp 1696145522
transform 1 0 3524 0 1 705
box -2 -3 26 103
use FILL  FILL_8_1
timestamp 1696145522
transform 1 0 3548 0 1 705
box -2 -3 10 103
use FILL  FILL_8_2
timestamp 1696145522
transform 1 0 3556 0 1 705
box -2 -3 10 103
use BUFX4  BUFX4_17
timestamp 1696145522
transform -1 0 36 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_196
timestamp 1696145522
transform -1 0 68 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_372
timestamp 1696145522
transform -1 0 92 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_227
timestamp 1696145522
transform 1 0 92 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_91
timestamp 1696145522
transform 1 0 116 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_41
timestamp 1696145522
transform -1 0 172 0 -1 905
box -2 -3 34 103
use INVX1  INVX1_38
timestamp 1696145522
transform -1 0 188 0 -1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_42
timestamp 1696145522
transform -1 0 220 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_274
timestamp 1696145522
transform -1 0 252 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_279
timestamp 1696145522
transform 1 0 252 0 -1 905
box -2 -3 26 103
use BUFX4  BUFX4_23
timestamp 1696145522
transform -1 0 308 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_340
timestamp 1696145522
transform -1 0 340 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_375
timestamp 1696145522
transform -1 0 372 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_109
timestamp 1696145522
transform -1 0 404 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_246
timestamp 1696145522
transform -1 0 428 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_411
timestamp 1696145522
transform -1 0 460 0 -1 905
box -2 -3 34 103
use INVX1  INVX1_104
timestamp 1696145522
transform 1 0 460 0 -1 905
box -2 -3 18 103
use FILL  FILL_8_0_0
timestamp 1696145522
transform -1 0 484 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_0_1
timestamp 1696145522
transform -1 0 492 0 -1 905
box -2 -3 10 103
use OAI21X1  OAI21X1_216
timestamp 1696145522
transform -1 0 524 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_411
timestamp 1696145522
transform -1 0 548 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_255
timestamp 1696145522
transform -1 0 580 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_385
timestamp 1696145522
transform -1 0 612 0 -1 905
box -2 -3 34 103
use INVX1  INVX1_60
timestamp 1696145522
transform -1 0 628 0 -1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_193
timestamp 1696145522
transform 1 0 628 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_39
timestamp 1696145522
transform -1 0 692 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_98
timestamp 1696145522
transform -1 0 724 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_596
timestamp 1696145522
transform -1 0 748 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_88
timestamp 1696145522
transform -1 0 772 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_99
timestamp 1696145522
transform -1 0 804 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_707
timestamp 1696145522
transform 1 0 804 0 -1 905
box -2 -3 34 103
use MUX2X1  MUX2X1_80
timestamp 1696145522
transform 1 0 836 0 -1 905
box -2 -3 50 103
use OAI21X1  OAI21X1_724
timestamp 1696145522
transform -1 0 916 0 -1 905
box -2 -3 34 103
use MUX2X1  MUX2X1_75
timestamp 1696145522
transform -1 0 964 0 -1 905
box -2 -3 50 103
use NAND2X1  NAND2X1_479
timestamp 1696145522
transform -1 0 988 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_295
timestamp 1696145522
transform -1 0 1012 0 -1 905
box -2 -3 26 103
use FILL  FILL_8_1_0
timestamp 1696145522
transform 1 0 1012 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_1_1
timestamp 1696145522
transform 1 0 1020 0 -1 905
box -2 -3 10 103
use AOI21X1  AOI21X1_329
timestamp 1696145522
transform 1 0 1028 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_763
timestamp 1696145522
transform 1 0 1060 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_796
timestamp 1696145522
transform -1 0 1124 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_245
timestamp 1696145522
transform -1 0 1148 0 -1 905
box -2 -3 26 103
use INVX1  INVX1_295
timestamp 1696145522
transform -1 0 1164 0 -1 905
box -2 -3 18 103
use NAND2X1  NAND2X1_447
timestamp 1696145522
transform -1 0 1188 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_555
timestamp 1696145522
transform 1 0 1188 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_330
timestamp 1696145522
transform 1 0 1220 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_128
timestamp 1696145522
transform -1 0 1276 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_848
timestamp 1696145522
transform -1 0 1308 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_815
timestamp 1696145522
transform 1 0 1308 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_816
timestamp 1696145522
transform 1 0 1340 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_785
timestamp 1696145522
transform -1 0 1404 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_213
timestamp 1696145522
transform -1 0 1428 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_817
timestamp 1696145522
transform -1 0 1460 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_694
timestamp 1696145522
transform -1 0 1492 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_170
timestamp 1696145522
transform -1 0 1516 0 -1 905
box -2 -3 26 103
use FILL  FILL_8_2_0
timestamp 1696145522
transform 1 0 1516 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_2_1
timestamp 1696145522
transform 1 0 1524 0 -1 905
box -2 -3 10 103
use OR2X2  OR2X2_10
timestamp 1696145522
transform 1 0 1532 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_808
timestamp 1696145522
transform -1 0 1596 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_461
timestamp 1696145522
transform 1 0 1596 0 -1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_462
timestamp 1696145522
transform 1 0 1620 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_829
timestamp 1696145522
transform 1 0 1644 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_636
timestamp 1696145522
transform -1 0 1700 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_728
timestamp 1696145522
transform 1 0 1700 0 -1 905
box -2 -3 34 103
use BUFX4  BUFX4_177
timestamp 1696145522
transform 1 0 1732 0 -1 905
box -2 -3 34 103
use BUFX4  BUFX4_186
timestamp 1696145522
transform 1 0 1764 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_830
timestamp 1696145522
transform 1 0 1796 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_800
timestamp 1696145522
transform -1 0 1860 0 -1 905
box -2 -3 34 103
use AND2X2  AND2X2_57
timestamp 1696145522
transform -1 0 1892 0 -1 905
box -2 -3 34 103
use BUFX4  BUFX4_115
timestamp 1696145522
transform 1 0 1892 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_789
timestamp 1696145522
transform -1 0 1956 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_235
timestamp 1696145522
transform 1 0 1956 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_786
timestamp 1696145522
transform -1 0 2012 0 -1 905
box -2 -3 34 103
use FILL  FILL_8_3_0
timestamp 1696145522
transform -1 0 2020 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_3_1
timestamp 1696145522
transform -1 0 2028 0 -1 905
box -2 -3 10 103
use OAI21X1  OAI21X1_695
timestamp 1696145522
transform -1 0 2060 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_810
timestamp 1696145522
transform 1 0 2060 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_809
timestamp 1696145522
transform -1 0 2124 0 -1 905
box -2 -3 34 103
use AOI22X1  AOI22X1_38
timestamp 1696145522
transform 1 0 2124 0 -1 905
box -2 -3 42 103
use AND2X2  AND2X2_62
timestamp 1696145522
transform 1 0 2164 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_797
timestamp 1696145522
transform 1 0 2196 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_698
timestamp 1696145522
transform 1 0 2228 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_300
timestamp 1696145522
transform -1 0 2292 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_227
timestamp 1696145522
transform -1 0 2316 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_850
timestamp 1696145522
transform 1 0 2316 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_849
timestamp 1696145522
transform 1 0 2348 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_342
timestamp 1696145522
transform 1 0 2380 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_619
timestamp 1696145522
transform -1 0 2436 0 -1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_341
timestamp 1696145522
transform 1 0 2436 0 -1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_66
timestamp 1696145522
transform -1 0 2500 0 -1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_348
timestamp 1696145522
transform 1 0 2500 0 -1 905
box -2 -3 34 103
use FILL  FILL_8_4_0
timestamp 1696145522
transform -1 0 2540 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_4_1
timestamp 1696145522
transform -1 0 2548 0 -1 905
box -2 -3 10 103
use BUFX4  BUFX4_2
timestamp 1696145522
transform -1 0 2580 0 -1 905
box -2 -3 34 103
use INVX4  INVX4_5
timestamp 1696145522
transform -1 0 2604 0 -1 905
box -2 -3 26 103
use CLKBUF1  CLKBUF1_7
timestamp 1696145522
transform -1 0 2676 0 -1 905
box -2 -3 74 103
use BUFX4  BUFX4_1
timestamp 1696145522
transform 1 0 2676 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_13
timestamp 1696145522
transform -1 0 2732 0 -1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_7
timestamp 1696145522
transform 1 0 2732 0 -1 905
box -2 -3 26 103
use INVX1  INVX1_5
timestamp 1696145522
transform -1 0 2772 0 -1 905
box -2 -3 18 103
use INVX2  INVX2_7
timestamp 1696145522
transform 1 0 2772 0 -1 905
box -2 -3 18 103
use NAND2X1  NAND2X1_16
timestamp 1696145522
transform 1 0 2788 0 -1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_13
timestamp 1696145522
transform 1 0 2812 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_18
timestamp 1696145522
transform -1 0 2860 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_865
timestamp 1696145522
transform 1 0 2860 0 -1 905
box -2 -3 34 103
use AND2X2  AND2X2_66
timestamp 1696145522
transform 1 0 2892 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_627
timestamp 1696145522
transform -1 0 2948 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_80
timestamp 1696145522
transform 1 0 2948 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_866
timestamp 1696145522
transform 1 0 2972 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_483
timestamp 1696145522
transform 1 0 3004 0 -1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_366
timestamp 1696145522
transform 1 0 3028 0 -1 905
box -2 -3 34 103
use FILL  FILL_8_5_0
timestamp 1696145522
transform 1 0 3060 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_5_1
timestamp 1696145522
transform 1 0 3068 0 -1 905
box -2 -3 10 103
use OAI21X1  OAI21X1_863
timestamp 1696145522
transform 1 0 3076 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_482
timestamp 1696145522
transform -1 0 3132 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_63
timestamp 1696145522
transform -1 0 3156 0 -1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_51
timestamp 1696145522
transform 1 0 3156 0 -1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_9
timestamp 1696145522
transform -1 0 3204 0 -1 905
box -2 -3 26 103
use INVX1  INVX1_7
timestamp 1696145522
transform -1 0 3220 0 -1 905
box -2 -3 18 103
use AND2X2  AND2X2_67
timestamp 1696145522
transform 1 0 3220 0 -1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_883
timestamp 1696145522
transform -1 0 3284 0 -1 905
box -2 -3 34 103
use XNOR2X1  XNOR2X1_15
timestamp 1696145522
transform -1 0 3340 0 -1 905
box -2 -3 58 103
use XOR2X1  XOR2X1_2
timestamp 1696145522
transform -1 0 3396 0 -1 905
box -2 -3 58 103
use BUFX4  BUFX4_15
timestamp 1696145522
transform -1 0 3428 0 -1 905
box -2 -3 34 103
use CLKBUF1  CLKBUF1_2
timestamp 1696145522
transform -1 0 3500 0 -1 905
box -2 -3 74 103
use BUFX2  BUFX2_19
timestamp 1696145522
transform 1 0 3500 0 -1 905
box -2 -3 26 103
use BUFX2  BUFX2_13
timestamp 1696145522
transform 1 0 3524 0 -1 905
box -2 -3 26 103
use FILL  FILL_9_1
timestamp 1696145522
transform -1 0 3556 0 -1 905
box -2 -3 10 103
use FILL  FILL_9_2
timestamp 1696145522
transform -1 0 3564 0 -1 905
box -2 -3 10 103
use NAND2X1  NAND2X1_229
timestamp 1696145522
transform -1 0 28 0 1 905
box -2 -3 26 103
use INVX1  INVX1_94
timestamp 1696145522
transform -1 0 44 0 1 905
box -2 -3 18 103
use INVX1  INVX1_113
timestamp 1696145522
transform 1 0 44 0 1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_256
timestamp 1696145522
transform 1 0 60 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_385
timestamp 1696145522
transform 1 0 92 0 1 905
box -2 -3 26 103
use INVX1  INVX1_114
timestamp 1696145522
transform 1 0 116 0 1 905
box -2 -3 18 103
use NAND2X1  NAND2X1_90
timestamp 1696145522
transform 1 0 132 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_399
timestamp 1696145522
transform -1 0 188 0 1 905
box -2 -3 34 103
use INVX1  INVX1_170
timestamp 1696145522
transform 1 0 188 0 1 905
box -2 -3 18 103
use NAND2X1  NAND2X1_352
timestamp 1696145522
transform -1 0 228 0 1 905
box -2 -3 26 103
use INVX1  INVX1_120
timestamp 1696145522
transform 1 0 228 0 1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_108
timestamp 1696145522
transform 1 0 244 0 1 905
box -2 -3 34 103
use INVX1  INVX1_62
timestamp 1696145522
transform -1 0 292 0 1 905
box -2 -3 18 103
use INVX1  INVX1_64
timestamp 1696145522
transform 1 0 292 0 1 905
box -2 -3 18 103
use NAND2X1  NAND2X1_390
timestamp 1696145522
transform -1 0 332 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_104
timestamp 1696145522
transform 1 0 332 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_154
timestamp 1696145522
transform 1 0 364 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_214
timestamp 1696145522
transform 1 0 388 0 1 905
box -2 -3 34 103
use MUX2X1  MUX2X1_26
timestamp 1696145522
transform 1 0 420 0 1 905
box -2 -3 50 103
use INVX1  INVX1_139
timestamp 1696145522
transform -1 0 484 0 1 905
box -2 -3 18 103
use FILL  FILL_9_0_0
timestamp 1696145522
transform 1 0 484 0 1 905
box -2 -3 10 103
use FILL  FILL_9_0_1
timestamp 1696145522
transform 1 0 492 0 1 905
box -2 -3 10 103
use INVX1  INVX1_150
timestamp 1696145522
transform 1 0 500 0 1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_321
timestamp 1696145522
transform 1 0 516 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_439
timestamp 1696145522
transform -1 0 580 0 1 905
box -2 -3 34 103
use INVX1  INVX1_124
timestamp 1696145522
transform 1 0 580 0 1 905
box -2 -3 18 103
use BUFX4  BUFX4_168
timestamp 1696145522
transform -1 0 628 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_341
timestamp 1696145522
transform -1 0 660 0 1 905
box -2 -3 34 103
use INVX1  INVX1_147
timestamp 1696145522
transform -1 0 676 0 1 905
box -2 -3 18 103
use NAND2X1  NAND2X1_143
timestamp 1696145522
transform 1 0 676 0 1 905
box -2 -3 26 103
use BUFX4  BUFX4_24
timestamp 1696145522
transform 1 0 700 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_748
timestamp 1696145522
transform -1 0 764 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_464
timestamp 1696145522
transform -1 0 788 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_144
timestamp 1696145522
transform 1 0 788 0 1 905
box -2 -3 26 103
use MUX2X1  MUX2X1_118
timestamp 1696145522
transform 1 0 812 0 1 905
box -2 -3 50 103
use NAND2X1  NAND2X1_569
timestamp 1696145522
transform 1 0 860 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_706
timestamp 1696145522
transform -1 0 916 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_727
timestamp 1696145522
transform 1 0 916 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_549
timestamp 1696145522
transform 1 0 948 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_485
timestamp 1696145522
transform 1 0 980 0 1 905
box -2 -3 34 103
use FILL  FILL_9_1_0
timestamp 1696145522
transform -1 0 1020 0 1 905
box -2 -3 10 103
use FILL  FILL_9_1_1
timestamp 1696145522
transform -1 0 1028 0 1 905
box -2 -3 10 103
use OAI21X1  OAI21X1_484
timestamp 1696145522
transform -1 0 1060 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_458
timestamp 1696145522
transform -1 0 1084 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_609
timestamp 1696145522
transform 1 0 1084 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_221
timestamp 1696145522
transform 1 0 1108 0 1 905
box -2 -3 34 103
use INVX8  INVX8_8
timestamp 1696145522
transform -1 0 1180 0 1 905
box -2 -3 42 103
use NOR2X1  NOR2X1_447
timestamp 1696145522
transform -1 0 1204 0 1 905
box -2 -3 26 103
use MUX2X1  MUX2X1_64
timestamp 1696145522
transform -1 0 1252 0 1 905
box -2 -3 50 103
use OAI22X1  OAI22X1_19
timestamp 1696145522
transform -1 0 1292 0 1 905
box -2 -3 42 103
use OAI22X1  OAI22X1_15
timestamp 1696145522
transform 1 0 1292 0 1 905
box -2 -3 42 103
use OAI21X1  OAI21X1_494
timestamp 1696145522
transform -1 0 1364 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_450
timestamp 1696145522
transform -1 0 1388 0 1 905
box -2 -3 26 103
use BUFX4  BUFX4_165
timestamp 1696145522
transform -1 0 1420 0 1 905
box -2 -3 34 103
use OAI22X1  OAI22X1_10
timestamp 1696145522
transform -1 0 1460 0 1 905
box -2 -3 42 103
use OAI21X1  OAI21X1_222
timestamp 1696145522
transform 1 0 1460 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_206
timestamp 1696145522
transform -1 0 1524 0 1 905
box -2 -3 34 103
use FILL  FILL_9_2_0
timestamp 1696145522
transform 1 0 1524 0 1 905
box -2 -3 10 103
use FILL  FILL_9_2_1
timestamp 1696145522
transform 1 0 1532 0 1 905
box -2 -3 10 103
use MUX2X1  MUX2X1_123
timestamp 1696145522
transform 1 0 1540 0 1 905
box -2 -3 50 103
use OAI21X1  OAI21X1_882
timestamp 1696145522
transform 1 0 1588 0 1 905
box -2 -3 34 103
use INVX8  INVX8_5
timestamp 1696145522
transform 1 0 1620 0 1 905
box -2 -3 42 103
use BUFX4  BUFX4_110
timestamp 1696145522
transform -1 0 1692 0 1 905
box -2 -3 34 103
use BUFX4  BUFX4_162
timestamp 1696145522
transform -1 0 1724 0 1 905
box -2 -3 34 103
use BUFX4  BUFX4_78
timestamp 1696145522
transform -1 0 1756 0 1 905
box -2 -3 34 103
use MUX2X1  MUX2X1_124
timestamp 1696145522
transform -1 0 1804 0 1 905
box -2 -3 50 103
use BUFX4  BUFX4_116
timestamp 1696145522
transform -1 0 1836 0 1 905
box -2 -3 34 103
use AND2X2  AND2X2_59
timestamp 1696145522
transform -1 0 1868 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_195
timestamp 1696145522
transform -1 0 1892 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_587
timestamp 1696145522
transform -1 0 1916 0 1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_427
timestamp 1696145522
transform -1 0 1940 0 1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_302
timestamp 1696145522
transform -1 0 1972 0 1 905
box -2 -3 34 103
use BUFX4  BUFX4_77
timestamp 1696145522
transform -1 0 2004 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_566
timestamp 1696145522
transform -1 0 2028 0 1 905
box -2 -3 26 103
use FILL  FILL_9_3_0
timestamp 1696145522
transform -1 0 2036 0 1 905
box -2 -3 10 103
use FILL  FILL_9_3_1
timestamp 1696145522
transform -1 0 2044 0 1 905
box -2 -3 10 103
use OAI22X1  OAI22X1_6
timestamp 1696145522
transform -1 0 2084 0 1 905
box -2 -3 42 103
use OAI21X1  OAI21X1_870
timestamp 1696145522
transform 1 0 2084 0 1 905
box -2 -3 34 103
use BUFX4  BUFX4_86
timestamp 1696145522
transform -1 0 2148 0 1 905
box -2 -3 34 103
use AND2X2  AND2X2_56
timestamp 1696145522
transform -1 0 2180 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_452
timestamp 1696145522
transform -1 0 2204 0 1 905
box -2 -3 26 103
use BUFX4  BUFX4_82
timestamp 1696145522
transform -1 0 2236 0 1 905
box -2 -3 34 103
use INVX1  INVX1_100
timestamp 1696145522
transform 1 0 2236 0 1 905
box -2 -3 18 103
use BUFX4  BUFX4_90
timestamp 1696145522
transform -1 0 2284 0 1 905
box -2 -3 34 103
use BUFX4  BUFX4_89
timestamp 1696145522
transform 1 0 2284 0 1 905
box -2 -3 34 103
use AND2X2  AND2X2_64
timestamp 1696145522
transform -1 0 2348 0 1 905
box -2 -3 34 103
use AND2X2  AND2X2_63
timestamp 1696145522
transform -1 0 2380 0 1 905
box -2 -3 34 103
use BUFX4  BUFX4_85
timestamp 1696145522
transform 1 0 2380 0 1 905
box -2 -3 34 103
use INVX8  INVX8_4
timestamp 1696145522
transform -1 0 2452 0 1 905
box -2 -3 42 103
use NAND2X1  NAND2X1_611
timestamp 1696145522
transform -1 0 2476 0 1 905
box -2 -3 26 103
use INVX2  INVX2_4
timestamp 1696145522
transform 1 0 2476 0 1 905
box -2 -3 18 103
use BUFX4  BUFX4_92
timestamp 1696145522
transform -1 0 2524 0 1 905
box -2 -3 34 103
use FILL  FILL_9_4_0
timestamp 1696145522
transform -1 0 2532 0 1 905
box -2 -3 10 103
use FILL  FILL_9_4_1
timestamp 1696145522
transform -1 0 2540 0 1 905
box -2 -3 10 103
use BUFX4  BUFX4_154
timestamp 1696145522
transform -1 0 2572 0 1 905
box -2 -3 34 103
use BUFX4  BUFX4_155
timestamp 1696145522
transform 1 0 2572 0 1 905
box -2 -3 34 103
use BUFX4  BUFX4_96
timestamp 1696145522
transform 1 0 2604 0 1 905
box -2 -3 34 103
use INVX4  INVX4_26
timestamp 1696145522
transform -1 0 2660 0 1 905
box -2 -3 26 103
use XNOR2X1  XNOR2X1_25
timestamp 1696145522
transform -1 0 2716 0 1 905
box -2 -3 58 103
use NOR2X1  NOR2X1_8
timestamp 1696145522
transform -1 0 2740 0 1 905
box -2 -3 26 103
use INVX1  INVX1_6
timestamp 1696145522
transform 1 0 2740 0 1 905
box -2 -3 18 103
use NAND2X1  NAND2X1_17
timestamp 1696145522
transform -1 0 2780 0 1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_49
timestamp 1696145522
transform -1 0 2804 0 1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_18
timestamp 1696145522
transform 1 0 2804 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_647
timestamp 1696145522
transform 1 0 2836 0 1 905
box -2 -3 34 103
use INVX1  INVX1_11
timestamp 1696145522
transform 1 0 2868 0 1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_7
timestamp 1696145522
transform 1 0 2884 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_19
timestamp 1696145522
transform -1 0 2940 0 1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_481
timestamp 1696145522
transform -1 0 2964 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_869
timestamp 1696145522
transform -1 0 2996 0 1 905
box -2 -3 34 103
use XNOR2X1  XNOR2X1_42
timestamp 1696145522
transform 1 0 2996 0 1 905
box -2 -3 58 103
use FILL  FILL_9_5_0
timestamp 1696145522
transform -1 0 3060 0 1 905
box -2 -3 10 103
use FILL  FILL_9_5_1
timestamp 1696145522
transform -1 0 3068 0 1 905
box -2 -3 10 103
use AOI21X1  AOI21X1_373
timestamp 1696145522
transform -1 0 3100 0 1 905
box -2 -3 34 103
use OR2X2  OR2X2_46
timestamp 1696145522
transform 1 0 3100 0 1 905
box -2 -3 34 103
use AOI21X1  AOI21X1_368
timestamp 1696145522
transform 1 0 3132 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_868
timestamp 1696145522
transform 1 0 3164 0 1 905
box -2 -3 34 103
use INVX2  INVX2_5
timestamp 1696145522
transform 1 0 3196 0 1 905
box -2 -3 18 103
use AOI22X1  AOI22X1_47
timestamp 1696145522
transform -1 0 3252 0 1 905
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_18
timestamp 1696145522
transform 1 0 3252 0 1 905
box -2 -3 98 103
use AOI22X1  AOI22X1_45
timestamp 1696145522
transform -1 0 3388 0 1 905
box -2 -3 42 103
use NAND3X1  NAND3X1_49
timestamp 1696145522
transform -1 0 3420 0 1 905
box -2 -3 34 103
use INVX1  INVX1_272
timestamp 1696145522
transform -1 0 3436 0 1 905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_17
timestamp 1696145522
transform 1 0 3436 0 1 905
box -2 -3 98 103
use BUFX2  BUFX2_20
timestamp 1696145522
transform 1 0 3532 0 1 905
box -2 -3 26 103
use FILL  FILL_10_1
timestamp 1696145522
transform 1 0 3556 0 1 905
box -2 -3 10 103
use OAI21X1  OAI21X1_292
timestamp 1696145522
transform -1 0 36 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_128
timestamp 1696145522
transform -1 0 52 0 -1 1105
box -2 -3 18 103
use INVX1  INVX1_42
timestamp 1696145522
transform 1 0 52 0 -1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_195
timestamp 1696145522
transform -1 0 100 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_93
timestamp 1696145522
transform -1 0 116 0 -1 1105
box -2 -3 18 103
use NAND2X1  NAND2X1_99
timestamp 1696145522
transform 1 0 116 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_339
timestamp 1696145522
transform 1 0 140 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_50
timestamp 1696145522
transform -1 0 204 0 -1 1105
box -2 -3 34 103
use BUFX4  BUFX4_19
timestamp 1696145522
transform 1 0 204 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_403
timestamp 1696145522
transform 1 0 236 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_431
timestamp 1696145522
transform -1 0 292 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_278
timestamp 1696145522
transform 1 0 292 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_301
timestamp 1696145522
transform -1 0 348 0 -1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_359
timestamp 1696145522
transform 1 0 348 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_351
timestamp 1696145522
transform 1 0 372 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_338
timestamp 1696145522
transform -1 0 428 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_325
timestamp 1696145522
transform -1 0 460 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_360
timestamp 1696145522
transform 1 0 460 0 -1 1105
box -2 -3 26 103
use FILL  FILL_10_0_0
timestamp 1696145522
transform -1 0 492 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_0_1
timestamp 1696145522
transform -1 0 500 0 -1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_353
timestamp 1696145522
transform -1 0 532 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_339
timestamp 1696145522
transform -1 0 556 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_326
timestamp 1696145522
transform -1 0 588 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_282
timestamp 1696145522
transform -1 0 620 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_351
timestamp 1696145522
transform 1 0 620 0 -1 1105
box -2 -3 26 103
use BUFX4  BUFX4_22
timestamp 1696145522
transform 1 0 644 0 -1 1105
box -2 -3 34 103
use MUX2X1  MUX2X1_27
timestamp 1696145522
transform 1 0 676 0 -1 1105
box -2 -3 50 103
use NAND2X1  NAND2X1_257
timestamp 1696145522
transform 1 0 724 0 -1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_621
timestamp 1696145522
transform 1 0 748 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_847
timestamp 1696145522
transform 1 0 772 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_761
timestamp 1696145522
transform 1 0 804 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_599
timestamp 1696145522
transform 1 0 836 0 -1 1105
box -2 -3 26 103
use INVX1  INVX1_299
timestamp 1696145522
transform 1 0 860 0 -1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_836
timestamp 1696145522
transform 1 0 876 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_261
timestamp 1696145522
transform -1 0 940 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_852
timestamp 1696145522
transform 1 0 940 0 -1 1105
box -2 -3 34 103
use AND2X2  AND2X2_61
timestamp 1696145522
transform 1 0 972 0 -1 1105
box -2 -3 34 103
use FILL  FILL_10_1_0
timestamp 1696145522
transform -1 0 1012 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_1_1
timestamp 1696145522
transform -1 0 1020 0 -1 1105
box -2 -3 10 103
use NAND2X1  NAND2X1_478
timestamp 1696145522
transform -1 0 1044 0 -1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_615
timestamp 1696145522
transform 1 0 1044 0 -1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_211
timestamp 1696145522
transform -1 0 1092 0 -1 1105
box -2 -3 26 103
use BUFX4  BUFX4_160
timestamp 1696145522
transform 1 0 1092 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_446
timestamp 1696145522
transform -1 0 1148 0 -1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_412
timestamp 1696145522
transform -1 0 1172 0 -1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_75
timestamp 1696145522
transform 1 0 1172 0 -1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_495
timestamp 1696145522
transform 1 0 1196 0 -1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_373
timestamp 1696145522
transform -1 0 1244 0 -1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_194
timestamp 1696145522
transform 1 0 1244 0 -1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_110
timestamp 1696145522
transform 1 0 1268 0 -1 1105
box -2 -3 26 103
use INVX1  INVX1_328
timestamp 1696145522
transform 1 0 1292 0 -1 1105
box -2 -3 18 103
use AOI21X1  AOI21X1_412
timestamp 1696145522
transform 1 0 1308 0 -1 1105
box -2 -3 34 103
use OAI22X1  OAI22X1_1
timestamp 1696145522
transform -1 0 1380 0 -1 1105
box -2 -3 42 103
use AOI21X1  AOI21X1_181
timestamp 1696145522
transform 1 0 1380 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_502
timestamp 1696145522
transform -1 0 1444 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_209
timestamp 1696145522
transform -1 0 1460 0 -1 1105
box -2 -3 18 103
use NOR2X1  NOR2X1_142
timestamp 1696145522
transform -1 0 1484 0 -1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_465
timestamp 1696145522
transform 1 0 1484 0 -1 1105
box -2 -3 26 103
use FILL  FILL_10_2_0
timestamp 1696145522
transform 1 0 1508 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_2_1
timestamp 1696145522
transform 1 0 1516 0 -1 1105
box -2 -3 10 103
use AOI21X1  AOI21X1_355
timestamp 1696145522
transform 1 0 1524 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_455
timestamp 1696145522
transform -1 0 1588 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_377
timestamp 1696145522
transform 1 0 1588 0 -1 1105
box -2 -3 34 103
use OAI22X1  OAI22X1_30
timestamp 1696145522
transform -1 0 1660 0 -1 1105
box -2 -3 42 103
use OAI21X1  OAI21X1_894
timestamp 1696145522
transform 1 0 1660 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_219
timestamp 1696145522
transform -1 0 1716 0 -1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_385
timestamp 1696145522
transform 1 0 1716 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_124
timestamp 1696145522
transform 1 0 1748 0 -1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_375
timestamp 1696145522
transform 1 0 1772 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_367
timestamp 1696145522
transform 1 0 1804 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_86
timestamp 1696145522
transform 1 0 1836 0 -1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_186
timestamp 1696145522
transform 1 0 1852 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_466
timestamp 1696145522
transform -1 0 1908 0 -1 1105
box -2 -3 26 103
use AND2X2  AND2X2_11
timestamp 1696145522
transform 1 0 1908 0 -1 1105
box -2 -3 34 103
use MUX2X1  MUX2X1_34
timestamp 1696145522
transform 1 0 1940 0 -1 1105
box -2 -3 50 103
use AOI21X1  AOI21X1_94
timestamp 1696145522
transform 1 0 1988 0 -1 1105
box -2 -3 34 103
use FILL  FILL_10_3_0
timestamp 1696145522
transform -1 0 2028 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_3_1
timestamp 1696145522
transform -1 0 2036 0 -1 1105
box -2 -3 10 103
use NOR2X1  NOR2X1_168
timestamp 1696145522
transform -1 0 2060 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_343
timestamp 1696145522
transform -1 0 2092 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_370
timestamp 1696145522
transform 1 0 2092 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_125
timestamp 1696145522
transform -1 0 2148 0 -1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_357
timestamp 1696145522
transform 1 0 2148 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_732
timestamp 1696145522
transform -1 0 2212 0 -1 1105
box -2 -3 34 103
use AND2X2  AND2X2_54
timestamp 1696145522
transform -1 0 2244 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_310
timestamp 1696145522
transform 1 0 2244 0 -1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_840
timestamp 1696145522
transform 1 0 2260 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_839
timestamp 1696145522
transform -1 0 2324 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_475
timestamp 1696145522
transform -1 0 2348 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_841
timestamp 1696145522
transform 1 0 2348 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_468
timestamp 1696145522
transform -1 0 2404 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_853
timestamp 1696145522
transform -1 0 2436 0 -1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_2
timestamp 1696145522
transform 1 0 2436 0 -1 1105
box -2 -3 98 103
use FILL  FILL_10_4_0
timestamp 1696145522
transform 1 0 2532 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_4_1
timestamp 1696145522
transform 1 0 2540 0 -1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_872
timestamp 1696145522
transform 1 0 2548 0 -1 1105
box -2 -3 34 103
use AND2X2  AND2X2_70
timestamp 1696145522
transform -1 0 2612 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_372
timestamp 1696145522
transform -1 0 2644 0 -1 1105
box -2 -3 34 103
use AOI22X1  AOI22X1_46
timestamp 1696145522
transform 1 0 2644 0 -1 1105
box -2 -3 42 103
use AOI21X1  AOI21X1_2
timestamp 1696145522
transform -1 0 2716 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_878
timestamp 1696145522
transform -1 0 2748 0 -1 1105
box -2 -3 34 103
use XNOR2X1  XNOR2X1_14
timestamp 1696145522
transform 1 0 2748 0 -1 1105
box -2 -3 58 103
use NAND2X1  NAND2X1_631
timestamp 1696145522
transform -1 0 2828 0 -1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_490
timestamp 1696145522
transform 1 0 2828 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_885
timestamp 1696145522
transform -1 0 2884 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_62
timestamp 1696145522
transform 1 0 2884 0 -1 1105
box -2 -3 26 103
use INVX1  INVX1_315
timestamp 1696145522
transform 1 0 2908 0 -1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_884
timestamp 1696145522
transform 1 0 2924 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_319
timestamp 1696145522
transform -1 0 2972 0 -1 1105
box -2 -3 18 103
use AOI21X1  AOI21X1_3
timestamp 1696145522
transform -1 0 3004 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_282
timestamp 1696145522
transform 1 0 3004 0 -1 1105
box -2 -3 18 103
use AOI21X1  AOI21X1_282
timestamp 1696145522
transform 1 0 3020 0 -1 1105
box -2 -3 34 103
use FILL  FILL_10_5_0
timestamp 1696145522
transform -1 0 3060 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_5_1
timestamp 1696145522
transform -1 0 3068 0 -1 1105
box -2 -3 10 103
use NOR2X1  NOR2X1_50
timestamp 1696145522
transform -1 0 3092 0 -1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_19
timestamp 1696145522
transform 1 0 3092 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_648
timestamp 1696145522
transform -1 0 3156 0 -1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_10
timestamp 1696145522
transform -1 0 3180 0 -1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_10
timestamp 1696145522
transform -1 0 3204 0 -1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_11
timestamp 1696145522
transform -1 0 3228 0 -1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_9
timestamp 1696145522
transform -1 0 3252 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_879
timestamp 1696145522
transform 1 0 3252 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_378
timestamp 1696145522
transform -1 0 3316 0 -1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_376
timestamp 1696145522
transform 1 0 3316 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_880
timestamp 1696145522
transform 1 0 3348 0 -1 1105
box -2 -3 34 103
use AOI22X1  AOI22X1_49
timestamp 1696145522
transform -1 0 3420 0 -1 1105
box -2 -3 42 103
use INVX1  INVX1_270
timestamp 1696145522
transform -1 0 3436 0 -1 1105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_20
timestamp 1696145522
transform 1 0 3436 0 -1 1105
box -2 -3 98 103
use BUFX2  BUFX2_22
timestamp 1696145522
transform 1 0 3532 0 -1 1105
box -2 -3 26 103
use FILL  FILL_11_1
timestamp 1696145522
transform -1 0 3564 0 -1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_201
timestamp 1696145522
transform 1 0 4 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_49
timestamp 1696145522
transform 1 0 36 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_40
timestamp 1696145522
transform -1 0 84 0 1 1105
box -2 -3 18 103
use NAND2X1  NAND2X1_280
timestamp 1696145522
transform -1 0 108 0 1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_228
timestamp 1696145522
transform 1 0 108 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_260
timestamp 1696145522
transform 1 0 132 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_350
timestamp 1696145522
transform -1 0 188 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_514
timestamp 1696145522
transform -1 0 220 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_296
timestamp 1696145522
transform -1 0 252 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_129
timestamp 1696145522
transform 1 0 252 0 1 1105
box -2 -3 18 103
use MUX2X1  MUX2X1_46
timestamp 1696145522
transform -1 0 316 0 1 1105
box -2 -3 50 103
use NAND2X1  NAND2X1_300
timestamp 1696145522
transform -1 0 340 0 1 1105
box -2 -3 26 103
use INVX1  INVX1_196
timestamp 1696145522
transform -1 0 356 0 1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_350
timestamp 1696145522
transform -1 0 388 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_277
timestamp 1696145522
transform 1 0 388 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_153
timestamp 1696145522
transform 1 0 420 0 1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_299
timestamp 1696145522
transform -1 0 468 0 1 1105
box -2 -3 26 103
use FILL  FILL_11_0_0
timestamp 1696145522
transform -1 0 476 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_0_1
timestamp 1696145522
transform -1 0 484 0 1 1105
box -2 -3 10 103
use MUX2X1  MUX2X1_49
timestamp 1696145522
transform -1 0 532 0 1 1105
box -2 -3 50 103
use NAND2X1  NAND2X1_334
timestamp 1696145522
transform 1 0 532 0 1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_300
timestamp 1696145522
transform -1 0 580 0 1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_284
timestamp 1696145522
transform -1 0 604 0 1 1105
box -2 -3 26 103
use MUX2X1  MUX2X1_25
timestamp 1696145522
transform -1 0 652 0 1 1105
box -2 -3 50 103
use OAI21X1  OAI21X1_40
timestamp 1696145522
transform -1 0 684 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_89
timestamp 1696145522
transform 1 0 684 0 1 1105
box -2 -3 26 103
use MUX2X1  MUX2X1_72
timestamp 1696145522
transform -1 0 756 0 1 1105
box -2 -3 50 103
use OAI21X1  OAI21X1_310
timestamp 1696145522
transform 1 0 756 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_327
timestamp 1696145522
transform -1 0 812 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_228
timestamp 1696145522
transform -1 0 844 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_678
timestamp 1696145522
transform 1 0 844 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_465
timestamp 1696145522
transform 1 0 876 0 1 1105
box -2 -3 26 103
use MUX2X1  MUX2X1_104
timestamp 1696145522
transform -1 0 948 0 1 1105
box -2 -3 50 103
use NAND2X1  NAND2X1_586
timestamp 1696145522
transform 1 0 948 0 1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_572
timestamp 1696145522
transform 1 0 972 0 1 1105
box -2 -3 26 103
use FILL  FILL_11_1_0
timestamp 1696145522
transform 1 0 996 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_1_1
timestamp 1696145522
transform 1 0 1004 0 1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_267
timestamp 1696145522
transform 1 0 1012 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_117
timestamp 1696145522
transform -1 0 1060 0 1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_826
timestamp 1696145522
transform -1 0 1092 0 1 1105
box -2 -3 34 103
use MUX2X1  MUX2X1_107
timestamp 1696145522
transform -1 0 1140 0 1 1105
box -2 -3 50 103
use MUX2X1  MUX2X1_105
timestamp 1696145522
transform -1 0 1188 0 1 1105
box -2 -3 50 103
use NAND2X1  NAND2X1_620
timestamp 1696145522
transform -1 0 1212 0 1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_274
timestamp 1696145522
transform -1 0 1236 0 1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_514
timestamp 1696145522
transform 1 0 1236 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_605
timestamp 1696145522
transform -1 0 1292 0 1 1105
box -2 -3 34 103
use MUX2X1  MUX2X1_122
timestamp 1696145522
transform 1 0 1292 0 1 1105
box -2 -3 50 103
use OAI21X1  OAI21X1_459
timestamp 1696145522
transform 1 0 1340 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_424
timestamp 1696145522
transform 1 0 1372 0 1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_449
timestamp 1696145522
transform -1 0 1420 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_123
timestamp 1696145522
transform -1 0 1452 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_570
timestamp 1696145522
transform -1 0 1484 0 1 1105
box -2 -3 34 103
use MUX2X1  MUX2X1_32
timestamp 1696145522
transform 1 0 1484 0 1 1105
box -2 -3 50 103
use FILL  FILL_11_2_0
timestamp 1696145522
transform 1 0 1532 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_2_1
timestamp 1696145522
transform 1 0 1540 0 1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_460
timestamp 1696145522
transform 1 0 1548 0 1 1105
box -2 -3 34 103
use MUX2X1  MUX2X1_127
timestamp 1696145522
transform 1 0 1580 0 1 1105
box -2 -3 50 103
use OAI21X1  OAI21X1_516
timestamp 1696145522
transform 1 0 1628 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_370
timestamp 1696145522
transform 1 0 1660 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_630
timestamp 1696145522
transform -1 0 1716 0 1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_145
timestamp 1696145522
transform 1 0 1716 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_860
timestamp 1696145522
transform 1 0 1740 0 1 1105
box -2 -3 34 103
use BUFX4  BUFX4_164
timestamp 1696145522
transform 1 0 1772 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_617
timestamp 1696145522
transform 1 0 1804 0 1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_428
timestamp 1696145522
transform -1 0 1852 0 1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_223
timestamp 1696145522
transform -1 0 1876 0 1 1105
box -2 -3 26 103
use INVX8  INVX8_9
timestamp 1696145522
transform 1 0 1876 0 1 1105
box -2 -3 42 103
use NOR2X1  NOR2X1_484
timestamp 1696145522
transform -1 0 1940 0 1 1105
box -2 -3 26 103
use OAI22X1  OAI22X1_28
timestamp 1696145522
transform -1 0 1980 0 1 1105
box -2 -3 42 103
use OAI21X1  OAI21X1_273
timestamp 1696145522
transform 1 0 1980 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_328
timestamp 1696145522
transform 1 0 2012 0 1 1105
box -2 -3 26 103
use FILL  FILL_11_3_0
timestamp 1696145522
transform 1 0 2036 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_3_1
timestamp 1696145522
transform 1 0 2044 0 1 1105
box -2 -3 10 103
use INVX1  INVX1_193
timestamp 1696145522
transform 1 0 2052 0 1 1105
box -2 -3 18 103
use AND2X2  AND2X2_69
timestamp 1696145522
transform 1 0 2068 0 1 1105
box -2 -3 34 103
use OR2X2  OR2X2_7
timestamp 1696145522
transform 1 0 2100 0 1 1105
box -2 -3 34 103
use BUFX4  BUFX4_84
timestamp 1696145522
transform 1 0 2132 0 1 1105
box -2 -3 34 103
use OAI22X1  OAI22X1_29
timestamp 1696145522
transform -1 0 2204 0 1 1105
box -2 -3 42 103
use AOI22X1  AOI22X1_7
timestamp 1696145522
transform -1 0 2244 0 1 1105
box -2 -3 42 103
use INVX8  INVX8_15
timestamp 1696145522
transform 1 0 2244 0 1 1105
box -2 -3 42 103
use OAI21X1  OAI21X1_203
timestamp 1696145522
transform 1 0 2284 0 1 1105
box -2 -3 34 103
use OR2X2  OR2X2_5
timestamp 1696145522
transform 1 0 2316 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_346
timestamp 1696145522
transform -1 0 2380 0 1 1105
box -2 -3 34 103
use BUFX4  BUFX4_87
timestamp 1696145522
transform 1 0 2380 0 1 1105
box -2 -3 34 103
use BUFX4  BUFX4_97
timestamp 1696145522
transform 1 0 2412 0 1 1105
box -2 -3 34 103
use AND2X2  AND2X2_53
timestamp 1696145522
transform 1 0 2444 0 1 1105
box -2 -3 34 103
use AOI22X1  AOI22X1_32
timestamp 1696145522
transform -1 0 2516 0 1 1105
box -2 -3 42 103
use AOI21X1  AOI21X1_74
timestamp 1696145522
transform 1 0 2516 0 1 1105
box -2 -3 34 103
use FILL  FILL_11_4_0
timestamp 1696145522
transform 1 0 2548 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_4_1
timestamp 1696145522
transform 1 0 2556 0 1 1105
box -2 -3 10 103
use INVX1  INVX1_268
timestamp 1696145522
transform 1 0 2564 0 1 1105
box -2 -3 18 103
use BUFX4  BUFX4_150
timestamp 1696145522
transform 1 0 2580 0 1 1105
box -2 -3 34 103
use BUFX4  BUFX4_152
timestamp 1696145522
transform 1 0 2612 0 1 1105
box -2 -3 34 103
use BUFX4  BUFX4_105
timestamp 1696145522
transform 1 0 2644 0 1 1105
box -2 -3 34 103
use BUFX4  BUFX4_100
timestamp 1696145522
transform 1 0 2676 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_364
timestamp 1696145522
transform 1 0 2708 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_629
timestamp 1696145522
transform -1 0 2764 0 1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_488
timestamp 1696145522
transform 1 0 2764 0 1 1105
box -2 -3 26 103
use AND2X2  AND2X2_68
timestamp 1696145522
transform 1 0 2788 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_876
timestamp 1696145522
transform 1 0 2820 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_877
timestamp 1696145522
transform -1 0 2884 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_317
timestamp 1696145522
transform -1 0 2900 0 1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_873
timestamp 1696145522
transform -1 0 2932 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_14
timestamp 1696145522
transform -1 0 2956 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_3
timestamp 1696145522
transform 1 0 2956 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_316
timestamp 1696145522
transform 1 0 2988 0 1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_26
timestamp 1696145522
transform 1 0 3004 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_66
timestamp 1696145522
transform 1 0 3036 0 1 1105
box -2 -3 26 103
use FILL  FILL_11_5_0
timestamp 1696145522
transform 1 0 3060 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_5_1
timestamp 1696145522
transform 1 0 3068 0 1 1105
box -2 -3 10 103
use NOR2X1  NOR2X1_485
timestamp 1696145522
transform 1 0 3076 0 1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_486
timestamp 1696145522
transform 1 0 3100 0 1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_12
timestamp 1696145522
transform 1 0 3124 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_874
timestamp 1696145522
transform 1 0 3148 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_489
timestamp 1696145522
transform -1 0 3204 0 1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_374
timestamp 1696145522
transform -1 0 3236 0 1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_881
timestamp 1696145522
transform 1 0 3236 0 1 1105
box -2 -3 34 103
use XNOR2X1  XNOR2X1_43
timestamp 1696145522
transform 1 0 3268 0 1 1105
box -2 -3 58 103
use BUFX2  BUFX2_4
timestamp 1696145522
transform 1 0 3324 0 1 1105
box -2 -3 26 103
use AOI22X1  AOI22X1_48
timestamp 1696145522
transform -1 0 3388 0 1 1105
box -2 -3 42 103
use NAND3X1  NAND3X1_48
timestamp 1696145522
transform -1 0 3420 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_271
timestamp 1696145522
transform -1 0 3436 0 1 1105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_19
timestamp 1696145522
transform 1 0 3436 0 1 1105
box -2 -3 98 103
use BUFX2  BUFX2_21
timestamp 1696145522
transform 1 0 3532 0 1 1105
box -2 -3 26 103
use FILL  FILL_12_1
timestamp 1696145522
transform 1 0 3556 0 1 1105
box -2 -3 10 103
use BUFX4  BUFX4_18
timestamp 1696145522
transform -1 0 36 0 -1 1305
box -2 -3 34 103
use MUX2X1  MUX2X1_42
timestamp 1696145522
transform -1 0 84 0 -1 1305
box -2 -3 50 103
use OAI21X1  OAI21X1_45
timestamp 1696145522
transform -1 0 116 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_39
timestamp 1696145522
transform -1 0 132 0 -1 1305
box -2 -3 18 103
use BUFX4  BUFX4_25
timestamp 1696145522
transform 1 0 132 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_187
timestamp 1696145522
transform 1 0 164 0 -1 1305
box -2 -3 18 103
use NAND2X1  NAND2X1_393
timestamp 1696145522
transform 1 0 180 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_458
timestamp 1696145522
transform 1 0 204 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_175
timestamp 1696145522
transform -1 0 252 0 -1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_415
timestamp 1696145522
transform -1 0 284 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_416
timestamp 1696145522
transform 1 0 284 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_537
timestamp 1696145522
transform 1 0 308 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_470
timestamp 1696145522
transform 1 0 340 0 -1 1305
box -2 -3 34 103
use BUFX4  BUFX4_122
timestamp 1696145522
transform 1 0 372 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_443
timestamp 1696145522
transform -1 0 436 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_331
timestamp 1696145522
transform 1 0 436 0 -1 1305
box -2 -3 26 103
use MUX2X1  MUX2X1_28
timestamp 1696145522
transform -1 0 508 0 -1 1305
box -2 -3 50 103
use FILL  FILL_12_0_0
timestamp 1696145522
transform -1 0 516 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_0_1
timestamp 1696145522
transform -1 0 524 0 -1 1305
box -2 -3 10 103
use BUFX4  BUFX4_166
timestamp 1696145522
transform -1 0 556 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_311
timestamp 1696145522
transform 1 0 556 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_419
timestamp 1696145522
transform 1 0 588 0 -1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_165
timestamp 1696145522
transform -1 0 636 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_446
timestamp 1696145522
transform -1 0 668 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_179
timestamp 1696145522
transform -1 0 700 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_183
timestamp 1696145522
transform -1 0 716 0 -1 1305
box -2 -3 18 103
use AOI21X1  AOI21X1_92
timestamp 1696145522
transform 1 0 716 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_135
timestamp 1696145522
transform 1 0 748 0 -1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_318
timestamp 1696145522
transform -1 0 796 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_234
timestamp 1696145522
transform -1 0 828 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_197
timestamp 1696145522
transform -1 0 852 0 -1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_381
timestamp 1696145522
transform -1 0 876 0 -1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_228
timestamp 1696145522
transform -1 0 900 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_185
timestamp 1696145522
transform -1 0 932 0 -1 1305
box -2 -3 34 103
use MUX2X1  MUX2X1_117
timestamp 1696145522
transform -1 0 980 0 -1 1305
box -2 -3 50 103
use NOR2X1  NOR2X1_287
timestamp 1696145522
transform -1 0 1004 0 -1 1305
box -2 -3 26 103
use FILL  FILL_12_1_0
timestamp 1696145522
transform -1 0 1012 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_1_1
timestamp 1696145522
transform -1 0 1020 0 -1 1305
box -2 -3 10 103
use NOR2X1  NOR2X1_294
timestamp 1696145522
transform -1 0 1044 0 -1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_212
timestamp 1696145522
transform 1 0 1044 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_416
timestamp 1696145522
transform 1 0 1068 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_361
timestamp 1696145522
transform -1 0 1124 0 -1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_148
timestamp 1696145522
transform 1 0 1124 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_417
timestamp 1696145522
transform 1 0 1156 0 -1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_382
timestamp 1696145522
transform 1 0 1180 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_119
timestamp 1696145522
transform 1 0 1212 0 -1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_376
timestamp 1696145522
transform -1 0 1260 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_204
timestamp 1696145522
transform 1 0 1260 0 -1 1305
box -2 -3 26 103
use OAI22X1  OAI22X1_16
timestamp 1696145522
transform -1 0 1324 0 -1 1305
box -2 -3 42 103
use OAI21X1  OAI21X1_945
timestamp 1696145522
transform -1 0 1356 0 -1 1305
box -2 -3 34 103
use AND2X2  AND2X2_25
timestamp 1696145522
transform 1 0 1356 0 -1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_40
timestamp 1696145522
transform 1 0 1388 0 -1 1305
box -2 -3 34 103
use AOI22X1  AOI22X1_58
timestamp 1696145522
transform -1 0 1460 0 -1 1305
box -2 -3 42 103
use INVX1  INVX1_261
timestamp 1696145522
transform 1 0 1460 0 -1 1305
box -2 -3 18 103
use NOR2X1  NOR2X1_368
timestamp 1696145522
transform -1 0 1500 0 -1 1305
box -2 -3 26 103
use FILL  FILL_12_2_0
timestamp 1696145522
transform -1 0 1508 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_2_1
timestamp 1696145522
transform -1 0 1516 0 -1 1305
box -2 -3 10 103
use OAI21X1  OAI21X1_524
timestamp 1696145522
transform -1 0 1548 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_468
timestamp 1696145522
transform -1 0 1572 0 -1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_160
timestamp 1696145522
transform -1 0 1596 0 -1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_420
timestamp 1696145522
transform 1 0 1596 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_449
timestamp 1696145522
transform -1 0 1652 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_377
timestamp 1696145522
transform 1 0 1652 0 -1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_135
timestamp 1696145522
transform -1 0 1716 0 -1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_78
timestamp 1696145522
transform 1 0 1716 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_494
timestamp 1696145522
transform 1 0 1748 0 -1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_457
timestamp 1696145522
transform -1 0 1796 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_515
timestamp 1696145522
transform -1 0 1828 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_474
timestamp 1696145522
transform 1 0 1828 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_538
timestamp 1696145522
transform -1 0 1884 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_637
timestamp 1696145522
transform -1 0 1908 0 -1 1305
box -2 -3 26 103
use OAI22X1  OAI22X1_31
timestamp 1696145522
transform 1 0 1908 0 -1 1305
box -2 -3 42 103
use NOR2X1  NOR2X1_493
timestamp 1696145522
transform -1 0 1972 0 -1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_187
timestamp 1696145522
transform -1 0 2004 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_296
timestamp 1696145522
transform -1 0 2028 0 -1 1305
box -2 -3 26 103
use FILL  FILL_12_3_0
timestamp 1696145522
transform -1 0 2036 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_3_1
timestamp 1696145522
transform -1 0 2044 0 -1 1305
box -2 -3 10 103
use AOI21X1  AOI21X1_196
timestamp 1696145522
transform -1 0 2076 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_221
timestamp 1696145522
transform -1 0 2092 0 -1 1305
box -2 -3 18 103
use AOI21X1  AOI21X1_120
timestamp 1696145522
transform -1 0 2124 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_313
timestamp 1696145522
transform 1 0 2124 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_867
timestamp 1696145522
transform -1 0 2188 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_442
timestamp 1696145522
transform -1 0 2212 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_237
timestamp 1696145522
transform 1 0 2212 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_448
timestamp 1696145522
transform 1 0 2244 0 -1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_264
timestamp 1696145522
transform -1 0 2292 0 -1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_149
timestamp 1696145522
transform -1 0 2324 0 -1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_93
timestamp 1696145522
transform 1 0 2324 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_340
timestamp 1696145522
transform 1 0 2356 0 -1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_63
timestamp 1696145522
transform 1 0 2380 0 -1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_66
timestamp 1696145522
transform 1 0 2412 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_435
timestamp 1696145522
transform -1 0 2468 0 -1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_146
timestamp 1696145522
transform -1 0 2492 0 -1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_172
timestamp 1696145522
transform 1 0 2492 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_305
timestamp 1696145522
transform 1 0 2524 0 -1 1305
box -2 -3 26 103
use FILL  FILL_12_4_0
timestamp 1696145522
transform -1 0 2556 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_4_1
timestamp 1696145522
transform -1 0 2564 0 -1 1305
box -2 -3 10 103
use NOR2X1  NOR2X1_149
timestamp 1696145522
transform -1 0 2588 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_699
timestamp 1696145522
transform -1 0 2620 0 -1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_47
timestamp 1696145522
transform 1 0 2620 0 -1 1305
box -2 -3 34 103
use INVX8  INVX8_14
timestamp 1696145522
transform 1 0 2652 0 -1 1305
box -2 -3 42 103
use BUFX4  BUFX4_3
timestamp 1696145522
transform -1 0 2724 0 -1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_69
timestamp 1696145522
transform 1 0 2724 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_633
timestamp 1696145522
transform 1 0 2756 0 -1 1305
box -2 -3 26 103
use AOI22X1  AOI22X1_51
timestamp 1696145522
transform -1 0 2820 0 -1 1305
box -2 -3 42 103
use INVX1  INVX1_321
timestamp 1696145522
transform -1 0 2836 0 -1 1305
box -2 -3 18 103
use NAND2X1  NAND2X1_638
timestamp 1696145522
transform -1 0 2860 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_897
timestamp 1696145522
transform -1 0 2892 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_495
timestamp 1696145522
transform 1 0 2892 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_4
timestamp 1696145522
transform 1 0 2916 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_14
timestamp 1696145522
transform -1 0 2972 0 -1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_6
timestamp 1696145522
transform 1 0 2972 0 -1 1305
box -2 -3 26 103
use INVX2  INVX2_3
timestamp 1696145522
transform -1 0 3012 0 -1 1305
box -2 -3 18 103
use NAND2X1  NAND2X1_632
timestamp 1696145522
transform -1 0 3036 0 -1 1305
box -2 -3 26 103
use FILL  FILL_12_5_0
timestamp 1696145522
transform -1 0 3044 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_5_1
timestamp 1696145522
transform -1 0 3052 0 -1 1305
box -2 -3 10 103
use XNOR2X1  XNOR2X1_13
timestamp 1696145522
transform -1 0 3108 0 -1 1305
box -2 -3 58 103
use NAND2X1  NAND2X1_7
timestamp 1696145522
transform 1 0 3108 0 -1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_52
timestamp 1696145522
transform -1 0 3156 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_649
timestamp 1696145522
transform 1 0 3156 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_8
timestamp 1696145522
transform -1 0 3212 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_650
timestamp 1696145522
transform -1 0 3244 0 -1 1305
box -2 -3 34 103
use BUFX4  BUFX4_12
timestamp 1696145522
transform -1 0 3276 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_628
timestamp 1696145522
transform 1 0 3276 0 -1 1305
box -2 -3 26 103
use OR2X2  OR2X2_47
timestamp 1696145522
transform 1 0 3300 0 -1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_70
timestamp 1696145522
transform -1 0 3364 0 -1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_890
timestamp 1696145522
transform 1 0 3364 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_635
timestamp 1696145522
transform -1 0 3420 0 -1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_403
timestamp 1696145522
transform 1 0 3420 0 -1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_401
timestamp 1696145522
transform -1 0 3468 0 -1 1305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_21
timestamp 1696145522
transform 1 0 3468 0 -1 1305
box -2 -3 98 103
use NAND2X1  NAND2X1_310
timestamp 1696145522
transform -1 0 28 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_234
timestamp 1696145522
transform -1 0 52 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_482
timestamp 1696145522
transform -1 0 84 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_98
timestamp 1696145522
transform 1 0 84 0 1 1305
box -2 -3 26 103
use BUFX4  BUFX4_120
timestamp 1696145522
transform 1 0 108 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_283
timestamp 1696145522
transform 1 0 140 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_456
timestamp 1696145522
transform 1 0 164 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_314
timestamp 1696145522
transform 1 0 188 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_423
timestamp 1696145522
transform 1 0 212 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_235
timestamp 1696145522
transform -1 0 268 0 1 1305
box -2 -3 34 103
use INVX1  INVX1_107
timestamp 1696145522
transform 1 0 268 0 1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_236
timestamp 1696145522
transform 1 0 284 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_233
timestamp 1696145522
transform 1 0 316 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_473
timestamp 1696145522
transform -1 0 372 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_431
timestamp 1696145522
transform 1 0 372 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_358
timestamp 1696145522
transform -1 0 420 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_483
timestamp 1696145522
transform -1 0 444 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_559
timestamp 1696145522
transform 1 0 444 0 1 1305
box -2 -3 34 103
use FILL  FILL_13_0_0
timestamp 1696145522
transform -1 0 484 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_0_1
timestamp 1696145522
transform -1 0 492 0 1 1305
box -2 -3 10 103
use OAI21X1  OAI21X1_506
timestamp 1696145522
transform -1 0 524 0 1 1305
box -2 -3 34 103
use MUX2X1  MUX2X1_44
timestamp 1696145522
transform 1 0 524 0 1 1305
box -2 -3 50 103
use NAND2X1  NAND2X1_329
timestamp 1696145522
transform -1 0 596 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_231
timestamp 1696145522
transform 1 0 596 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_260
timestamp 1696145522
transform 1 0 628 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_212
timestamp 1696145522
transform 1 0 652 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_365
timestamp 1696145522
transform 1 0 676 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_308
timestamp 1696145522
transform 1 0 708 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_366
timestamp 1696145522
transform 1 0 740 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_261
timestamp 1696145522
transform 1 0 764 0 1 1305
box -2 -3 26 103
use MUX2X1  MUX2X1_29
timestamp 1696145522
transform 1 0 788 0 1 1305
box -2 -3 50 103
use INVX1  INVX1_167
timestamp 1696145522
transform 1 0 836 0 1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_390
timestamp 1696145522
transform 1 0 852 0 1 1305
box -2 -3 34 103
use INVX1  INVX1_168
timestamp 1696145522
transform 1 0 884 0 1 1305
box -2 -3 18 103
use NAND2X1  NAND2X1_218
timestamp 1696145522
transform -1 0 924 0 1 1305
box -2 -3 26 103
use BUFX4  BUFX4_21
timestamp 1696145522
transform 1 0 924 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_558
timestamp 1696145522
transform 1 0 956 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_269
timestamp 1696145522
transform -1 0 1012 0 1 1305
box -2 -3 34 103
use FILL  FILL_13_1_0
timestamp 1696145522
transform -1 0 1020 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_1_1
timestamp 1696145522
transform -1 0 1028 0 1 1305
box -2 -3 10 103
use NAND2X1  NAND2X1_291
timestamp 1696145522
transform -1 0 1052 0 1 1305
box -2 -3 26 103
use MUX2X1  MUX2X1_39
timestamp 1696145522
transform 1 0 1052 0 1 1305
box -2 -3 50 103
use AOI21X1  AOI21X1_354
timestamp 1696145522
transform 1 0 1100 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_150
timestamp 1696145522
transform -1 0 1156 0 1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_79
timestamp 1696145522
transform -1 0 1188 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_301
timestamp 1696145522
transform 1 0 1188 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_560
timestamp 1696145522
transform 1 0 1212 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_299
timestamp 1696145522
transform -1 0 1268 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_561
timestamp 1696145522
transform 1 0 1268 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_391
timestamp 1696145522
transform 1 0 1300 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_497
timestamp 1696145522
transform -1 0 1356 0 1 1305
box -2 -3 26 103
use MUX2X1  MUX2X1_126
timestamp 1696145522
transform 1 0 1356 0 1 1305
box -2 -3 50 103
use OAI21X1  OAI21X1_403
timestamp 1696145522
transform 1 0 1404 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_404
timestamp 1696145522
transform 1 0 1436 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_398
timestamp 1696145522
transform 1 0 1468 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_367
timestamp 1696145522
transform -1 0 1524 0 1 1305
box -2 -3 26 103
use FILL  FILL_13_2_0
timestamp 1696145522
transform -1 0 1532 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_2_1
timestamp 1696145522
transform -1 0 1540 0 1 1305
box -2 -3 10 103
use NAND2X1  NAND2X1_623
timestamp 1696145522
transform -1 0 1564 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_539
timestamp 1696145522
transform -1 0 1596 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_193
timestamp 1696145522
transform -1 0 1620 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_386
timestamp 1696145522
transform 1 0 1620 0 1 1305
box -2 -3 34 103
use MUX2X1  MUX2X1_128
timestamp 1696145522
transform 1 0 1652 0 1 1305
box -2 -3 50 103
use BUFX4  BUFX4_79
timestamp 1696145522
transform -1 0 1732 0 1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_20
timestamp 1696145522
transform 1 0 1732 0 1 1305
box -2 -3 34 103
use BUFX4  BUFX4_163
timestamp 1696145522
transform 1 0 1764 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_887
timestamp 1696145522
transform 1 0 1796 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_395
timestamp 1696145522
transform -1 0 1852 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_420
timestamp 1696145522
transform 1 0 1852 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_396
timestamp 1696145522
transform -1 0 1908 0 1 1305
box -2 -3 26 103
use AOI22X1  AOI22X1_12
timestamp 1696145522
transform -1 0 1948 0 1 1305
box -2 -3 42 103
use AND2X2  AND2X2_18
timestamp 1696145522
transform 1 0 1948 0 1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_122
timestamp 1696145522
transform 1 0 1980 0 1 1305
box -2 -3 34 103
use FILL  FILL_13_3_0
timestamp 1696145522
transform -1 0 2020 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_3_1
timestamp 1696145522
transform -1 0 2028 0 1 1305
box -2 -3 10 103
use AOI21X1  AOI21X1_121
timestamp 1696145522
transform -1 0 2060 0 1 1305
box -2 -3 34 103
use AOI22X1  AOI22X1_50
timestamp 1696145522
transform -1 0 2100 0 1 1305
box -2 -3 42 103
use NAND3X1  NAND3X1_18
timestamp 1696145522
transform 1 0 2100 0 1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_362
timestamp 1696145522
transform -1 0 2164 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_355
timestamp 1696145522
transform 1 0 2164 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_448
timestamp 1696145522
transform 1 0 2196 0 1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_105
timestamp 1696145522
transform 1 0 2228 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_483
timestamp 1696145522
transform 1 0 2260 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_253
timestamp 1696145522
transform -1 0 2316 0 1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_252
timestamp 1696145522
transform -1 0 2340 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_317
timestamp 1696145522
transform -1 0 2372 0 1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_168
timestamp 1696145522
transform -1 0 2404 0 1 1305
box -2 -3 34 103
use INVX4  INVX4_11
timestamp 1696145522
transform 1 0 2404 0 1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_196
timestamp 1696145522
transform -1 0 2452 0 1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_199
timestamp 1696145522
transform 1 0 2452 0 1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_198
timestamp 1696145522
transform -1 0 2500 0 1 1305
box -2 -3 26 103
use NAND3X1  NAND3X1_24
timestamp 1696145522
transform 1 0 2500 0 1 1305
box -2 -3 34 103
use FILL  FILL_13_4_0
timestamp 1696145522
transform -1 0 2540 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_4_1
timestamp 1696145522
transform -1 0 2548 0 1 1305
box -2 -3 10 103
use OAI21X1  OAI21X1_496
timestamp 1696145522
transform -1 0 2580 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_271
timestamp 1696145522
transform 1 0 2580 0 1 1305
box -2 -3 34 103
use AOI22X1  AOI22X1_15
timestamp 1696145522
transform -1 0 2652 0 1 1305
box -2 -3 42 103
use OAI21X1  OAI21X1_490
timestamp 1696145522
transform 1 0 2652 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_497
timestamp 1696145522
transform -1 0 2716 0 1 1305
box -2 -3 34 103
use AOI22X1  AOI22X1_19
timestamp 1696145522
transform -1 0 2756 0 1 1305
box -2 -3 42 103
use OAI21X1  OAI21X1_871
timestamp 1696145522
transform 1 0 2756 0 1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_371
timestamp 1696145522
transform -1 0 2820 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_889
timestamp 1696145522
transform 1 0 2820 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_132
timestamp 1696145522
transform 1 0 2852 0 1 1305
box -2 -3 26 103
use BUFX4  BUFX4_173
timestamp 1696145522
transform 1 0 2876 0 1 1305
box -2 -3 34 103
use AND2X2  AND2X2_52
timestamp 1696145522
transform -1 0 2940 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_861
timestamp 1696145522
transform 1 0 2940 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_862
timestamp 1696145522
transform -1 0 3004 0 1 1305
box -2 -3 34 103
use BUFX4  BUFX4_91
timestamp 1696145522
transform -1 0 3036 0 1 1305
box -2 -3 34 103
use FILL  FILL_13_5_0
timestamp 1696145522
transform -1 0 3044 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_5_1
timestamp 1696145522
transform -1 0 3052 0 1 1305
box -2 -3 10 103
use BUFX4  BUFX4_140
timestamp 1696145522
transform -1 0 3084 0 1 1305
box -2 -3 34 103
use BUFX4  BUFX4_108
timestamp 1696145522
transform 1 0 3084 0 1 1305
box -2 -3 34 103
use XNOR2X1  XNOR2X1_12
timestamp 1696145522
transform 1 0 3116 0 1 1305
box -2 -3 58 103
use OAI21X1  OAI21X1_896
timestamp 1696145522
transform 1 0 3172 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_895
timestamp 1696145522
transform -1 0 3236 0 1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_491
timestamp 1696145522
transform -1 0 3260 0 1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_492
timestamp 1696145522
transform 1 0 3260 0 1 1305
box -2 -3 26 103
use BUFX4  BUFX4_138
timestamp 1696145522
transform 1 0 3284 0 1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_386
timestamp 1696145522
transform -1 0 3348 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_893
timestamp 1696145522
transform -1 0 3380 0 1 1305
box -2 -3 34 103
use XNOR2X1  XNOR2X1_45
timestamp 1696145522
transform -1 0 3436 0 1 1305
box -2 -3 58 103
use OAI21X1  OAI21X1_5
timestamp 1696145522
transform -1 0 3468 0 1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_381
timestamp 1696145522
transform 1 0 3468 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_886
timestamp 1696145522
transform 1 0 3500 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_634
timestamp 1696145522
transform -1 0 3556 0 1 1305
box -2 -3 26 103
use FILL  FILL_14_1
timestamp 1696145522
transform 1 0 3556 0 1 1305
box -2 -3 10 103
use INVX1  INVX1_96
timestamp 1696145522
transform 1 0 4 0 -1 1505
box -2 -3 18 103
use OAI21X1  OAI21X1_200
timestamp 1696145522
transform 1 0 20 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_374
timestamp 1696145522
transform 1 0 52 0 -1 1505
box -2 -3 34 103
use INVX1  INVX1_160
timestamp 1696145522
transform -1 0 100 0 -1 1505
box -2 -3 18 103
use NAND2X1  NAND2X1_371
timestamp 1696145522
transform 1 0 100 0 -1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_282
timestamp 1696145522
transform 1 0 124 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_259
timestamp 1696145522
transform -1 0 180 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_338
timestamp 1696145522
transform -1 0 212 0 -1 1505
box -2 -3 34 103
use MUX2X1  MUX2X1_38
timestamp 1696145522
transform -1 0 260 0 -1 1505
box -2 -3 50 103
use OAI21X1  OAI21X1_414
timestamp 1696145522
transform -1 0 292 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_266
timestamp 1696145522
transform 1 0 292 0 -1 1505
box -2 -3 26 103
use INVX1  INVX1_181
timestamp 1696145522
transform -1 0 332 0 -1 1505
box -2 -3 18 103
use NOR2X1  NOR2X1_266
timestamp 1696145522
transform -1 0 356 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_505
timestamp 1696145522
transform -1 0 388 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_631
timestamp 1696145522
transform 1 0 388 0 -1 1505
box -2 -3 34 103
use OAI22X1  OAI22X1_23
timestamp 1696145522
transform 1 0 420 0 -1 1505
box -2 -3 42 103
use OAI21X1  OAI21X1_324
timestamp 1696145522
transform -1 0 492 0 -1 1505
box -2 -3 34 103
use FILL  FILL_14_0_0
timestamp 1696145522
transform -1 0 500 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_0_1
timestamp 1696145522
transform -1 0 508 0 -1 1505
box -2 -3 10 103
use MUX2X1  MUX2X1_43
timestamp 1696145522
transform -1 0 556 0 -1 1505
box -2 -3 50 103
use MUX2X1  MUX2X1_37
timestamp 1696145522
transform -1 0 604 0 -1 1505
box -2 -3 50 103
use OAI21X1  OAI21X1_220
timestamp 1696145522
transform 1 0 604 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_251
timestamp 1696145522
transform -1 0 660 0 -1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_365
timestamp 1696145522
transform 1 0 660 0 -1 1505
box -2 -3 26 103
use BUFX4  BUFX4_16
timestamp 1696145522
transform 1 0 684 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_325
timestamp 1696145522
transform 1 0 716 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_225
timestamp 1696145522
transform 1 0 740 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_346
timestamp 1696145522
transform 1 0 772 0 -1 1505
box -2 -3 26 103
use INVX1  INVX1_146
timestamp 1696145522
transform 1 0 796 0 -1 1505
box -2 -3 18 103
use OAI21X1  OAI21X1_332
timestamp 1696145522
transform 1 0 812 0 -1 1505
box -2 -3 34 103
use INVX1  INVX1_134
timestamp 1696145522
transform 1 0 844 0 -1 1505
box -2 -3 18 103
use OAI21X1  OAI21X1_309
timestamp 1696145522
transform 1 0 860 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_326
timestamp 1696145522
transform -1 0 916 0 -1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_136
timestamp 1696145522
transform 1 0 916 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_247
timestamp 1696145522
transform 1 0 940 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_271
timestamp 1696145522
transform 1 0 972 0 -1 1505
box -2 -3 26 103
use FILL  FILL_14_1_0
timestamp 1696145522
transform 1 0 996 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_1_1
timestamp 1696145522
transform 1 0 1004 0 -1 1505
box -2 -3 10 103
use MUX2X1  MUX2X1_120
timestamp 1696145522
transform 1 0 1012 0 -1 1505
box -2 -3 50 103
use MUX2X1  MUX2X1_111
timestamp 1696145522
transform -1 0 1108 0 -1 1505
box -2 -3 50 103
use MUX2X1  MUX2X1_112
timestamp 1696145522
transform -1 0 1156 0 -1 1505
box -2 -3 50 103
use OAI21X1  OAI21X1_85
timestamp 1696145522
transform -1 0 1188 0 -1 1505
box -2 -3 34 103
use AND2X2  AND2X2_23
timestamp 1696145522
transform 1 0 1188 0 -1 1505
box -2 -3 34 103
use AND2X2  AND2X2_20
timestamp 1696145522
transform 1 0 1220 0 -1 1505
box -2 -3 34 103
use BUFX4  BUFX4_167
timestamp 1696145522
transform 1 0 1252 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_645
timestamp 1696145522
transform -1 0 1308 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_784
timestamp 1696145522
transform 1 0 1308 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_615
timestamp 1696145522
transform 1 0 1340 0 -1 1505
box -2 -3 34 103
use MUX2X1  MUX2X1_116
timestamp 1696145522
transform 1 0 1372 0 -1 1505
box -2 -3 50 103
use MUX2X1  MUX2X1_125
timestamp 1696145522
transform 1 0 1420 0 -1 1505
box -2 -3 50 103
use NAND2X1  NAND2X1_508
timestamp 1696145522
transform -1 0 1492 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_908
timestamp 1696145522
transform 1 0 1492 0 -1 1505
box -2 -3 34 103
use FILL  FILL_14_2_0
timestamp 1696145522
transform -1 0 1532 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_2_1
timestamp 1696145522
transform -1 0 1540 0 -1 1505
box -2 -3 10 103
use INVX2  INVX2_48
timestamp 1696145522
transform -1 0 1556 0 -1 1505
box -2 -3 18 103
use AOI21X1  AOI21X1_391
timestamp 1696145522
transform 1 0 1556 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_498
timestamp 1696145522
transform -1 0 1612 0 -1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_388
timestamp 1696145522
transform 1 0 1612 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_81
timestamp 1696145522
transform -1 0 1668 0 -1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_396
timestamp 1696145522
transform 1 0 1668 0 -1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_406
timestamp 1696145522
transform 1 0 1700 0 -1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_315
timestamp 1696145522
transform 1 0 1732 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_502
timestamp 1696145522
transform -1 0 1788 0 -1 1505
box -2 -3 26 103
use INVX1  INVX1_320
timestamp 1696145522
transform 1 0 1788 0 -1 1505
box -2 -3 18 103
use OAI21X1  OAI21X1_625
timestamp 1696145522
transform 1 0 1804 0 -1 1505
box -2 -3 34 103
use OAI22X1  OAI22X1_21
timestamp 1696145522
transform 1 0 1836 0 -1 1505
box -2 -3 42 103
use NAND2X1  NAND2X1_520
timestamp 1696145522
transform 1 0 1876 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_419
timestamp 1696145522
transform 1 0 1900 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_366
timestamp 1696145522
transform -1 0 1964 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_80
timestamp 1696145522
transform -1 0 1988 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_616
timestamp 1696145522
transform -1 0 2020 0 -1 1505
box -2 -3 34 103
use FILL  FILL_14_3_0
timestamp 1696145522
transform -1 0 2028 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_3_1
timestamp 1696145522
transform -1 0 2036 0 -1 1505
box -2 -3 10 103
use BUFX4  BUFX4_81
timestamp 1696145522
transform -1 0 2068 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_497
timestamp 1696145522
transform -1 0 2092 0 -1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_116
timestamp 1696145522
transform -1 0 2124 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_447
timestamp 1696145522
transform 1 0 2124 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_87
timestamp 1696145522
transform 1 0 2156 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_875
timestamp 1696145522
transform -1 0 2212 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_471
timestamp 1696145522
transform 1 0 2212 0 -1 1505
box -2 -3 34 103
use BUFX4  BUFX4_161
timestamp 1696145522
transform -1 0 2276 0 -1 1505
box -2 -3 34 103
use BUFX4  BUFX4_159
timestamp 1696145522
transform -1 0 2308 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_268
timestamp 1696145522
transform 1 0 2308 0 -1 1505
box -2 -3 26 103
use BUFX4  BUFX4_170
timestamp 1696145522
transform -1 0 2364 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_487
timestamp 1696145522
transform 1 0 2364 0 -1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_180
timestamp 1696145522
transform -1 0 2420 0 -1 1505
box -2 -3 34 103
use OAI22X1  OAI22X1_8
timestamp 1696145522
transform -1 0 2460 0 -1 1505
box -2 -3 42 103
use NAND2X1  NAND2X1_276
timestamp 1696145522
transform -1 0 2484 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_466
timestamp 1696145522
transform 1 0 2484 0 -1 1505
box -2 -3 34 103
use INVX1  INVX1_195
timestamp 1696145522
transform 1 0 2516 0 -1 1505
box -2 -3 18 103
use FILL  FILL_14_4_0
timestamp 1696145522
transform -1 0 2540 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_4_1
timestamp 1696145522
transform -1 0 2548 0 -1 1505
box -2 -3 10 103
use INVX1  INVX1_189
timestamp 1696145522
transform -1 0 2564 0 -1 1505
box -2 -3 18 103
use AOI21X1  AOI21X1_155
timestamp 1696145522
transform 1 0 2564 0 -1 1505
box -2 -3 34 103
use AND2X2  AND2X2_14
timestamp 1696145522
transform 1 0 2596 0 -1 1505
box -2 -3 34 103
use BUFX4  BUFX4_172
timestamp 1696145522
transform 1 0 2628 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_272
timestamp 1696145522
transform -1 0 2684 0 -1 1505
box -2 -3 26 103
use INVX1  INVX1_110
timestamp 1696145522
transform 1 0 2684 0 -1 1505
box -2 -3 18 103
use OAI21X1  OAI21X1_252
timestamp 1696145522
transform 1 0 2700 0 -1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_72
timestamp 1696145522
transform 1 0 2732 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_715
timestamp 1696145522
transform -1 0 2796 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_431
timestamp 1696145522
transform 1 0 2796 0 -1 1505
box -2 -3 26 103
use INVX1  INVX1_111
timestamp 1696145522
transform 1 0 2820 0 -1 1505
box -2 -3 18 103
use OAI21X1  OAI21X1_262
timestamp 1696145522
transform -1 0 2868 0 -1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_75
timestamp 1696145522
transform -1 0 2900 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_473
timestamp 1696145522
transform 1 0 2900 0 -1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_477
timestamp 1696145522
transform -1 0 2948 0 -1 1505
box -2 -3 26 103
use AOI22X1  AOI22X1_31
timestamp 1696145522
transform -1 0 2988 0 -1 1505
box -2 -3 42 103
use NAND2X1  NAND2X1_265
timestamp 1696145522
transform -1 0 3012 0 -1 1505
box -2 -3 26 103
use INVX1  INVX1_269
timestamp 1696145522
transform -1 0 3028 0 -1 1505
box -2 -3 18 103
use AOI21X1  AOI21X1_379
timestamp 1696145522
transform 1 0 3028 0 -1 1505
box -2 -3 34 103
use FILL  FILL_14_5_0
timestamp 1696145522
transform 1 0 3060 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_5_1
timestamp 1696145522
transform 1 0 3068 0 -1 1505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_1
timestamp 1696145522
transform 1 0 3076 0 -1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_892
timestamp 1696145522
transform -1 0 3204 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_891
timestamp 1696145522
transform -1 0 3236 0 -1 1505
box -2 -3 34 103
use AND2X2  AND2X2_71
timestamp 1696145522
transform 1 0 3236 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_898
timestamp 1696145522
transform -1 0 3300 0 -1 1505
box -2 -3 34 103
use AND2X2  AND2X2_72
timestamp 1696145522
transform -1 0 3332 0 -1 1505
box -2 -3 34 103
use OR2X2  OR2X2_48
timestamp 1696145522
transform -1 0 3364 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_61
timestamp 1696145522
transform 1 0 3364 0 -1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_283
timestamp 1696145522
transform -1 0 3420 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_2
timestamp 1696145522
transform -1 0 3452 0 -1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_5
timestamp 1696145522
transform -1 0 3476 0 -1 1505
box -2 -3 26 103
use BUFX4  BUFX4_13
timestamp 1696145522
transform -1 0 3508 0 -1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_20
timestamp 1696145522
transform -1 0 3540 0 -1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_5
timestamp 1696145522
transform -1 0 3564 0 -1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_558
timestamp 1696145522
transform -1 0 84 0 -1 1705
box -2 -3 34 103
use MUX2X1  MUX2X1_58
timestamp 1696145522
transform -1 0 52 0 -1 1705
box -2 -3 50 103
use NAND2X1  NAND2X1_233
timestamp 1696145522
transform 1 0 36 0 1 1505
box -2 -3 26 103
use BUFX4  BUFX4_126
timestamp 1696145522
transform -1 0 36 0 1 1505
box -2 -3 34 103
use BUFX4  BUFX4_69
timestamp 1696145522
transform 1 0 108 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_370
timestamp 1696145522
transform 1 0 84 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_373
timestamp 1696145522
transform -1 0 116 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_441
timestamp 1696145522
transform 1 0 60 0 1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_263
timestamp 1696145522
transform 1 0 140 0 -1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_313
timestamp 1696145522
transform -1 0 172 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_295
timestamp 1696145522
transform 1 0 116 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_406
timestamp 1696145522
transform 1 0 164 0 -1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_349
timestamp 1696145522
transform 1 0 172 0 1 1505
box -2 -3 26 103
use MUX2X1  MUX2X1_47
timestamp 1696145522
transform 1 0 220 0 -1 1705
box -2 -3 50 103
use OAI21X1  OAI21X1_434
timestamp 1696145522
transform -1 0 220 0 -1 1705
box -2 -3 34 103
use MUX2X1  MUX2X1_40
timestamp 1696145522
transform 1 0 196 0 1 1505
box -2 -3 50 103
use OAI21X1  OAI21X1_402
timestamp 1696145522
transform -1 0 300 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_392
timestamp 1696145522
transform -1 0 292 0 1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_373
timestamp 1696145522
transform -1 0 268 0 1 1505
box -2 -3 26 103
use MUX2X1  MUX2X1_52
timestamp 1696145522
transform -1 0 380 0 -1 1705
box -2 -3 50 103
use OAI21X1  OAI21X1_578
timestamp 1696145522
transform 1 0 300 0 -1 1705
box -2 -3 34 103
use MUX2X1  MUX2X1_63
timestamp 1696145522
transform 1 0 324 0 1 1505
box -2 -3 50 103
use OAI21X1  OAI21X1_469
timestamp 1696145522
transform 1 0 292 0 1 1505
box -2 -3 34 103
use MUX2X1  MUX2X1_67
timestamp 1696145522
transform 1 0 380 0 -1 1705
box -2 -3 50 103
use OAI21X1  OAI21X1_442
timestamp 1696145522
transform -1 0 428 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_267
timestamp 1696145522
transform 1 0 372 0 1 1505
box -2 -3 26 103
use MUX2X1  MUX2X1_55
timestamp 1696145522
transform 1 0 428 0 -1 1705
box -2 -3 50 103
use NAND2X1  NAND2X1_337
timestamp 1696145522
transform 1 0 452 0 1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_415
timestamp 1696145522
transform 1 0 428 0 1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_273
timestamp 1696145522
transform 1 0 524 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_493
timestamp 1696145522
transform 1 0 492 0 -1 1705
box -2 -3 34 103
use FILL  FILL_16_0_1
timestamp 1696145522
transform 1 0 484 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_0_0
timestamp 1696145522
transform 1 0 476 0 -1 1705
box -2 -3 10 103
use NAND2X1  NAND2X1_379
timestamp 1696145522
transform -1 0 548 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_384
timestamp 1696145522
transform 1 0 492 0 1 1505
box -2 -3 34 103
use FILL  FILL_15_0_1
timestamp 1696145522
transform 1 0 484 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_0_0
timestamp 1696145522
transform 1 0 476 0 1 1505
box -2 -3 10 103
use NOR2X1  NOR2X1_139
timestamp 1696145522
transform -1 0 604 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_66
timestamp 1696145522
transform 1 0 548 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_312
timestamp 1696145522
transform 1 0 572 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_100
timestamp 1696145522
transform -1 0 572 0 1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_71
timestamp 1696145522
transform 1 0 620 0 -1 1705
box -2 -3 34 103
use INVX1  INVX1_106
timestamp 1696145522
transform -1 0 620 0 -1 1705
box -2 -3 18 103
use OAI21X1  OAI21X1_87
timestamp 1696145522
transform 1 0 604 0 1 1505
box -2 -3 34 103
use INVX1  INVX1_109
timestamp 1696145522
transform 1 0 652 0 -1 1705
box -2 -3 18 103
use OAI21X1  OAI21X1_88
timestamp 1696145522
transform -1 0 668 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_178
timestamp 1696145522
transform 1 0 684 0 -1 1705
box -2 -3 34 103
use INVX1  INVX1_52
timestamp 1696145522
transform -1 0 684 0 -1 1705
box -2 -3 18 103
use INVX1  INVX1_53
timestamp 1696145522
transform 1 0 692 0 1 1505
box -2 -3 18 103
use NOR2X1  NOR2X1_83
timestamp 1696145522
transform -1 0 692 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_248
timestamp 1696145522
transform -1 0 748 0 -1 1705
box -2 -3 34 103
use BUFX4  BUFX4_124
timestamp 1696145522
transform 1 0 724 0 1 1505
box -2 -3 34 103
use INVX1  INVX1_55
timestamp 1696145522
transform 1 0 708 0 1 1505
box -2 -3 18 103
use OAI21X1  OAI21X1_128
timestamp 1696145522
transform 1 0 748 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_117
timestamp 1696145522
transform 1 0 756 0 1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_169
timestamp 1696145522
transform -1 0 804 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_74
timestamp 1696145522
transform -1 0 812 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_405
timestamp 1696145522
transform -1 0 860 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_388
timestamp 1696145522
transform 1 0 804 0 -1 1705
box -2 -3 26 103
use OR2X2  OR2X2_13
timestamp 1696145522
transform 1 0 836 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_254
timestamp 1696145522
transform 1 0 812 0 1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_274
timestamp 1696145522
transform -1 0 884 0 -1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_293
timestamp 1696145522
transform 1 0 868 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_426
timestamp 1696145522
transform 1 0 900 0 -1 1705
box -2 -3 34 103
use INVX1  INVX1_88
timestamp 1696145522
transform 1 0 884 0 -1 1705
box -2 -3 18 103
use OAI21X1  OAI21X1_268
timestamp 1696145522
transform -1 0 940 0 1 1505
box -2 -3 34 103
use INVX1  INVX1_73
timestamp 1696145522
transform 1 0 892 0 1 1505
box -2 -3 18 103
use OAI21X1  OAI21X1_265
timestamp 1696145522
transform 1 0 956 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_182
timestamp 1696145522
transform 1 0 932 0 -1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_101
timestamp 1696145522
transform -1 0 964 0 1 1505
box -2 -3 26 103
use MUX2X1  MUX2X1_33
timestamp 1696145522
transform -1 0 1052 0 -1 1705
box -2 -3 50 103
use FILL  FILL_16_1_1
timestamp 1696145522
transform -1 0 1004 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_1_0
timestamp 1696145522
transform -1 0 996 0 -1 1705
box -2 -3 10 103
use FILL  FILL_15_1_0
timestamp 1696145522
transform 1 0 1012 0 1 1505
box -2 -3 10 103
use NAND2X1  NAND2X1_397
timestamp 1696145522
transform -1 0 1012 0 1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_294
timestamp 1696145522
transform 1 0 964 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_139
timestamp 1696145522
transform -1 0 1084 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_726
timestamp 1696145522
transform -1 0 1092 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_272
timestamp 1696145522
transform 1 0 1028 0 1 1505
box -2 -3 34 103
use FILL  FILL_15_1_1
timestamp 1696145522
transform 1 0 1020 0 1 1505
box -2 -3 10 103
use INVX1  INVX1_118
timestamp 1696145522
transform -1 0 1100 0 -1 1705
box -2 -3 18 103
use OAI21X1  OAI21X1_79
timestamp 1696145522
transform 1 0 1140 0 -1 1705
box -2 -3 34 103
use INVX1  INVX1_293
timestamp 1696145522
transform -1 0 1140 0 -1 1705
box -2 -3 18 103
use NOR2X1  NOR2X1_151
timestamp 1696145522
transform -1 0 1124 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_134
timestamp 1696145522
transform -1 0 1172 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_172
timestamp 1696145522
transform 1 0 1116 0 1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_585
timestamp 1696145522
transform -1 0 1116 0 1 1505
box -2 -3 26 103
use MUX2X1  MUX2X1_121
timestamp 1696145522
transform -1 0 1220 0 -1 1705
box -2 -3 50 103
use OAI21X1  OAI21X1_145
timestamp 1696145522
transform 1 0 1172 0 1 1505
box -2 -3 34 103
use MUX2X1  MUX2X1_36
timestamp 1696145522
transform 1 0 1220 0 -1 1705
box -2 -3 50 103
use OAI21X1  OAI21X1_342
timestamp 1696145522
transform 1 0 1228 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_188
timestamp 1696145522
transform 1 0 1204 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_251
timestamp 1696145522
transform 1 0 1268 0 -1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_84
timestamp 1696145522
transform -1 0 1284 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_250
timestamp 1696145522
transform -1 0 1332 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_734
timestamp 1696145522
transform -1 0 1316 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_548
timestamp 1696145522
transform -1 0 1364 0 -1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_360
timestamp 1696145522
transform -1 0 1364 0 1 1505
box -2 -3 26 103
use NAND2X1  NAND2X1_605
timestamp 1696145522
transform 1 0 1316 0 1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_204
timestamp 1696145522
transform 1 0 1364 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_333
timestamp 1696145522
transform -1 0 1396 0 1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_227
timestamp 1696145522
transform 1 0 1396 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_513
timestamp 1696145522
transform -1 0 1420 0 1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_206
timestamp 1696145522
transform -1 0 1452 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_356
timestamp 1696145522
transform 1 0 1420 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_406
timestamp 1696145522
transform 1 0 1476 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_519
timestamp 1696145522
transform -1 0 1476 0 -1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_177
timestamp 1696145522
transform -1 0 1508 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_89
timestamp 1696145522
transform 1 0 1452 0 1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_241
timestamp 1696145522
transform -1 0 1556 0 -1 1705
box -2 -3 34 103
use FILL  FILL_16_2_1
timestamp 1696145522
transform -1 0 1524 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_2_0
timestamp 1696145522
transform -1 0 1516 0 -1 1705
box -2 -3 10 103
use NAND2X1  NAND2X1_643
timestamp 1696145522
transform -1 0 1548 0 1 1505
box -2 -3 26 103
use FILL  FILL_15_2_1
timestamp 1696145522
transform -1 0 1524 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_2_0
timestamp 1696145522
transform -1 0 1516 0 1 1505
box -2 -3 10 103
use AOI21X1  AOI21X1_243
timestamp 1696145522
transform 1 0 1556 0 -1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_144
timestamp 1696145522
transform -1 0 1580 0 1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_228
timestamp 1696145522
transform 1 0 1588 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_435
timestamp 1696145522
transform -1 0 1612 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_925
timestamp 1696145522
transform -1 0 1652 0 -1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_107
timestamp 1696145522
transform 1 0 1612 0 1 1505
box -2 -3 34 103
use OAI22X1  OAI22X1_32
timestamp 1696145522
transform -1 0 1708 0 -1 1705
box -2 -3 42 103
use INVX1  INVX1_324
timestamp 1696145522
transform -1 0 1668 0 -1 1705
box -2 -3 18 103
use NOR2X1  NOR2X1_176
timestamp 1696145522
transform 1 0 1676 0 1 1505
box -2 -3 26 103
use AND2X2  AND2X2_7
timestamp 1696145522
transform 1 0 1644 0 1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_409
timestamp 1696145522
transform -1 0 1764 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_480
timestamp 1696145522
transform -1 0 1732 0 -1 1705
box -2 -3 26 103
use OAI22X1  OAI22X1_33
timestamp 1696145522
transform -1 0 1740 0 1 1505
box -2 -3 42 103
use MUX2X1  MUX2X1_129
timestamp 1696145522
transform 1 0 1764 0 -1 1705
box -2 -3 50 103
use AOI21X1  AOI21X1_108
timestamp 1696145522
transform -1 0 1804 0 1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_106
timestamp 1696145522
transform 1 0 1740 0 1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_404
timestamp 1696145522
transform 1 0 1812 0 -1 1705
box -2 -3 34 103
use INVX1  INVX1_151
timestamp 1696145522
transform -1 0 1820 0 1 1505
box -2 -3 18 103
use OAI22X1  OAI22X1_18
timestamp 1696145522
transform 1 0 1844 0 -1 1705
box -2 -3 42 103
use OAI22X1  OAI22X1_14
timestamp 1696145522
transform 1 0 1820 0 1 1505
box -2 -3 42 103
use OAI21X1  OAI21X1_933
timestamp 1696145522
transform 1 0 1884 0 -1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_242
timestamp 1696145522
transform 1 0 1892 0 1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_212
timestamp 1696145522
transform 1 0 1860 0 1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_220
timestamp 1696145522
transform 1 0 1940 0 -1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_205
timestamp 1696145522
transform -1 0 1940 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_562
timestamp 1696145522
transform -1 0 1972 0 1 1505
box -2 -3 34 103
use INVX1  INVX1_228
timestamp 1696145522
transform -1 0 1940 0 1 1505
box -2 -3 18 103
use OAI22X1  OAI22X1_37
timestamp 1696145522
transform -1 0 2012 0 -1 1705
box -2 -3 42 103
use NOR2X1  NOR2X1_317
timestamp 1696145522
transform -1 0 1996 0 1 1505
box -2 -3 26 103
use FILL  FILL_16_3_1
timestamp 1696145522
transform -1 0 2052 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_3_0
timestamp 1696145522
transform -1 0 2044 0 -1 1705
box -2 -3 10 103
use NOR2X1  NOR2X1_502
timestamp 1696145522
transform 1 0 2012 0 -1 1705
box -2 -3 26 103
use MUX2X1  MUX2X1_48
timestamp 1696145522
transform -1 0 2092 0 1 1505
box -2 -3 50 103
use FILL  FILL_15_3_1
timestamp 1696145522
transform -1 0 2044 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_3_0
timestamp 1696145522
transform -1 0 2036 0 1 1505
box -2 -3 10 103
use OAI21X1  OAI21X1_528
timestamp 1696145522
transform -1 0 2028 0 1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_226
timestamp 1696145522
transform -1 0 2116 0 -1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_400
timestamp 1696145522
transform -1 0 2084 0 -1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_268
timestamp 1696145522
transform -1 0 2124 0 1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_127
timestamp 1696145522
transform -1 0 2180 0 -1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_128
timestamp 1696145522
transform 1 0 2116 0 -1 1705
box -2 -3 34 103
use MUX2X1  MUX2X1_21
timestamp 1696145522
transform 1 0 2124 0 1 1505
box -2 -3 50 103
use NAND2X1  NAND2X1_125
timestamp 1696145522
transform 1 0 2172 0 1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_36
timestamp 1696145522
transform 1 0 2212 0 -1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_86
timestamp 1696145522
transform 1 0 2180 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_86
timestamp 1696145522
transform -1 0 2228 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_90
timestamp 1696145522
transform 1 0 2244 0 -1 1705
box -2 -3 34 103
use INVX1  INVX1_54
timestamp 1696145522
transform 1 0 2244 0 1 1505
box -2 -3 18 103
use INVX2  INVX2_49
timestamp 1696145522
transform 1 0 2228 0 1 1505
box -2 -3 18 103
use AOI21X1  AOI21X1_41
timestamp 1696145522
transform -1 0 2308 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_507
timestamp 1696145522
transform -1 0 2292 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_189
timestamp 1696145522
transform 1 0 2308 0 -1 1705
box -2 -3 26 103
use OR2X2  OR2X2_31
timestamp 1696145522
transform 1 0 2316 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_477
timestamp 1696145522
transform 1 0 2292 0 1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_203
timestamp 1696145522
transform -1 0 2364 0 -1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_183
timestamp 1696145522
transform -1 0 2380 0 1 1505
box -2 -3 34 103
use OAI22X1  OAI22X1_2
timestamp 1696145522
transform -1 0 2404 0 -1 1705
box -2 -3 42 103
use OAI21X1  OAI21X1_508
timestamp 1696145522
transform -1 0 2412 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_318
timestamp 1696145522
transform -1 0 2460 0 -1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_91
timestamp 1696145522
transform -1 0 2436 0 -1 1705
box -2 -3 34 103
use INVX1  INVX1_56
timestamp 1696145522
transform -1 0 2452 0 1 1505
box -2 -3 18 103
use NAND2X1  NAND2X1_452
timestamp 1696145522
transform -1 0 2436 0 1 1505
box -2 -3 26 103
use OAI22X1  OAI22X1_27
timestamp 1696145522
transform 1 0 2460 0 -1 1705
box -2 -3 42 103
use NAND3X1  NAND3X1_15
timestamp 1696145522
transform -1 0 2516 0 1 1505
box -2 -3 34 103
use OR2X2  OR2X2_16
timestamp 1696145522
transform 1 0 2452 0 1 1505
box -2 -3 34 103
use FILL  FILL_16_4_0
timestamp 1696145522
transform 1 0 2532 0 -1 1705
box -2 -3 10 103
use OAI21X1  OAI21X1_749
timestamp 1696145522
transform 1 0 2500 0 -1 1705
box -2 -3 34 103
use OR2X2  OR2X2_15
timestamp 1696145522
transform 1 0 2516 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_523
timestamp 1696145522
transform 1 0 2548 0 -1 1705
box -2 -3 34 103
use FILL  FILL_16_4_1
timestamp 1696145522
transform 1 0 2540 0 -1 1705
box -2 -3 10 103
use AOI21X1  AOI21X1_100
timestamp 1696145522
transform 1 0 2564 0 1 1505
box -2 -3 34 103
use FILL  FILL_15_4_1
timestamp 1696145522
transform 1 0 2556 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_4_0
timestamp 1696145522
transform 1 0 2548 0 1 1505
box -2 -3 10 103
use NAND2X1  NAND2X1_286
timestamp 1696145522
transform -1 0 2628 0 -1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_140
timestamp 1696145522
transform -1 0 2604 0 -1 1705
box -2 -3 26 103
use AOI21X1  AOI21X1_101
timestamp 1696145522
transform 1 0 2596 0 1 1505
box -2 -3 34 103
use BUFX4  BUFX4_176
timestamp 1696145522
transform -1 0 2660 0 -1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_235
timestamp 1696145522
transform -1 0 2652 0 1 1505
box -2 -3 26 103
use AND2X2  AND2X2_22
timestamp 1696145522
transform 1 0 2684 0 -1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_402
timestamp 1696145522
transform -1 0 2684 0 -1 1705
box -2 -3 26 103
use AOI21X1  AOI21X1_160
timestamp 1696145522
transform 1 0 2684 0 1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_154
timestamp 1696145522
transform 1 0 2652 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_813
timestamp 1696145522
transform 1 0 2716 0 -1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_239
timestamp 1696145522
transform -1 0 2740 0 1 1505
box -2 -3 26 103
use BUFX4  BUFX4_80
timestamp 1696145522
transform -1 0 2780 0 -1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_25
timestamp 1696145522
transform 1 0 2740 0 1 1505
box -2 -3 34 103
use BUFX4  BUFX4_9
timestamp 1696145522
transform -1 0 2812 0 -1 1705
box -2 -3 34 103
use OR2X2  OR2X2_27
timestamp 1696145522
transform -1 0 2804 0 1 1505
box -2 -3 34 103
use BUFX4  BUFX4_10
timestamp 1696145522
transform -1 0 2844 0 -1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_161
timestamp 1696145522
transform -1 0 2836 0 1 1505
box -2 -3 34 103
use BUFX4  BUFX4_7
timestamp 1696145522
transform 1 0 2844 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_465
timestamp 1696145522
transform -1 0 2868 0 1 1505
box -2 -3 34 103
use BUFX4  BUFX4_175
timestamp 1696145522
transform 1 0 2876 0 -1 1705
box -2 -3 34 103
use OR2X2  OR2X2_25
timestamp 1696145522
transform -1 0 2924 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_129
timestamp 1696145522
transform -1 0 2892 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_436
timestamp 1696145522
transform -1 0 2940 0 -1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_67
timestamp 1696145522
transform -1 0 2956 0 1 1505
box -2 -3 34 103
use OR2X2  OR2X2_44
timestamp 1696145522
transform 1 0 2972 0 -1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_143
timestamp 1696145522
transform 1 0 2940 0 -1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_467
timestamp 1696145522
transform -1 0 2980 0 1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_89
timestamp 1696145522
transform 1 0 3004 0 -1 1705
box -2 -3 26 103
use NAND3X1  NAND3X1_8
timestamp 1696145522
transform 1 0 2980 0 1 1505
box -2 -3 34 103
use FILL  FILL_16_5_0
timestamp 1696145522
transform 1 0 3044 0 -1 1705
box -2 -3 10 103
use INVX1  INVX1_57
timestamp 1696145522
transform -1 0 3044 0 -1 1705
box -2 -3 18 103
use FILL  FILL_15_5_1
timestamp 1696145522
transform 1 0 3044 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_5_0
timestamp 1696145522
transform 1 0 3036 0 1 1505
box -2 -3 10 103
use NOR2X1  NOR2X1_478
timestamp 1696145522
transform -1 0 3036 0 1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_77
timestamp 1696145522
transform 1 0 3060 0 -1 1705
box -2 -3 26 103
use FILL  FILL_16_5_1
timestamp 1696145522
transform 1 0 3052 0 -1 1705
box -2 -3 10 103
use BUFX4  BUFX4_65
timestamp 1696145522
transform 1 0 3052 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_90
timestamp 1696145522
transform -1 0 3180 0 -1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_79
timestamp 1696145522
transform -1 0 3156 0 -1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_88
timestamp 1696145522
transform 1 0 3108 0 -1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_86
timestamp 1696145522
transform -1 0 3108 0 -1 1705
box -2 -3 26 103
use NAND3X1  NAND3X1_71
timestamp 1696145522
transform -1 0 3180 0 1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_392
timestamp 1696145522
transform 1 0 3116 0 1 1505
box -2 -3 34 103
use BUFX4  BUFX4_83
timestamp 1696145522
transform 1 0 3084 0 1 1505
box -2 -3 34 103
use AOI22X1  AOI22X1_53
timestamp 1696145522
transform 1 0 3252 0 -1 1705
box -2 -3 42 103
use BUFX4  BUFX4_60
timestamp 1696145522
transform -1 0 3252 0 -1 1705
box -2 -3 34 103
use INVX1  INVX1_51
timestamp 1696145522
transform -1 0 3220 0 -1 1705
box -2 -3 18 103
use NAND2X1  NAND2X1_640
timestamp 1696145522
transform -1 0 3204 0 -1 1705
box -2 -3 26 103
use AOI21X1  AOI21X1_380
timestamp 1696145522
transform 1 0 3204 0 1 1505
box -2 -3 34 103
use INVX4  INVX4_3
timestamp 1696145522
transform 1 0 3180 0 1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_22
timestamp 1696145522
transform 1 0 3236 0 1 1505
box -2 -3 98 103
use AOI21X1  AOI21X1_4
timestamp 1696145522
transform 1 0 3292 0 -1 1705
box -2 -3 34 103
use INVX1  INVX1_8
timestamp 1696145522
transform 1 0 3324 0 -1 1705
box -2 -3 18 103
use AND2X2  AND2X2_73
timestamp 1696145522
transform -1 0 3364 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_15
timestamp 1696145522
transform -1 0 3388 0 -1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_11
timestamp 1696145522
transform -1 0 3364 0 -1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_496
timestamp 1696145522
transform -1 0 3388 0 1 1505
box -2 -3 26 103
use OAI21X1  OAI21X1_6
timestamp 1696145522
transform -1 0 3420 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_900
timestamp 1696145522
transform -1 0 3420 0 1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_5
timestamp 1696145522
transform 1 0 3420 0 -1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_899
timestamp 1696145522
transform -1 0 3452 0 1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_27
timestamp 1696145522
transform 1 0 3476 0 -1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_6
timestamp 1696145522
transform 1 0 3452 0 -1 1705
box -2 -3 26 103
use AOI21X1  AOI21X1_384
timestamp 1696145522
transform -1 0 3484 0 1 1505
box -2 -3 34 103
use NAND2X1  NAND2X1_66
timestamp 1696145522
transform -1 0 3532 0 -1 1705
box -2 -3 26 103
use AOI21X1  AOI21X1_389
timestamp 1696145522
transform -1 0 3540 0 1 1505
box -2 -3 34 103
use BUFX2  BUFX2_3
timestamp 1696145522
transform 1 0 3484 0 1 1505
box -2 -3 26 103
use FILL  FILL_17_1
timestamp 1696145522
transform -1 0 3556 0 -1 1705
box -2 -3 10 103
use INVX1  INVX1_28
timestamp 1696145522
transform 1 0 3532 0 -1 1705
box -2 -3 18 103
use NAND2X1  NAND2X1_536
timestamp 1696145522
transform -1 0 3564 0 1 1505
box -2 -3 26 103
use FILL  FILL_17_2
timestamp 1696145522
transform -1 0 3564 0 -1 1705
box -2 -3 10 103
use OAI21X1  OAI21X1_593
timestamp 1696145522
transform -1 0 36 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_510
timestamp 1696145522
transform -1 0 60 0 1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_482
timestamp 1696145522
transform -1 0 84 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_630
timestamp 1696145522
transform 1 0 84 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_94
timestamp 1696145522
transform 1 0 116 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_125
timestamp 1696145522
transform -1 0 172 0 1 1705
box -2 -3 34 103
use BUFX4  BUFX4_121
timestamp 1696145522
transform 1 0 172 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_629
timestamp 1696145522
transform -1 0 236 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_387
timestamp 1696145522
transform 1 0 236 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_481
timestamp 1696145522
transform 1 0 260 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_430
timestamp 1696145522
transform 1 0 292 0 1 1705
box -2 -3 26 103
use INVX2  INVX2_57
timestamp 1696145522
transform -1 0 332 0 1 1705
box -2 -3 18 103
use NOR2X1  NOR2X1_99
timestamp 1696145522
transform 1 0 332 0 1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_501
timestamp 1696145522
transform -1 0 380 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_536
timestamp 1696145522
transform -1 0 412 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_568
timestamp 1696145522
transform -1 0 444 0 1 1705
box -2 -3 34 103
use MUX2X1  MUX2X1_54
timestamp 1696145522
transform 1 0 444 0 1 1705
box -2 -3 50 103
use FILL  FILL_17_0_0
timestamp 1696145522
transform 1 0 492 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_0_1
timestamp 1696145522
transform 1 0 500 0 1 1705
box -2 -3 10 103
use NAND2X1  NAND2X1_446
timestamp 1696145522
transform 1 0 508 0 1 1705
box -2 -3 26 103
use AOI21X1  AOI21X1_235
timestamp 1696145522
transform 1 0 532 0 1 1705
box -2 -3 34 103
use AOI22X1  AOI22X1_26
timestamp 1696145522
transform 1 0 564 0 1 1705
box -2 -3 42 103
use NAND2X1  NAND2X1_149
timestamp 1696145522
transform 1 0 604 0 1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_113
timestamp 1696145522
transform -1 0 652 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_249
timestamp 1696145522
transform 1 0 652 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_275
timestamp 1696145522
transform -1 0 708 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_301
timestamp 1696145522
transform 1 0 708 0 1 1705
box -2 -3 34 103
use BUFX4  BUFX4_118
timestamp 1696145522
transform 1 0 740 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_73
timestamp 1696145522
transform 1 0 772 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_211
timestamp 1696145522
transform -1 0 828 0 1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_316
timestamp 1696145522
transform -1 0 852 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_299
timestamp 1696145522
transform -1 0 884 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_184
timestamp 1696145522
transform 1 0 884 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_401
timestamp 1696145522
transform -1 0 940 0 1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_321
timestamp 1696145522
transform 1 0 940 0 1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_290
timestamp 1696145522
transform 1 0 964 0 1 1705
box -2 -3 26 103
use FILL  FILL_17_1_0
timestamp 1696145522
transform 1 0 988 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_1_1
timestamp 1696145522
transform 1 0 996 0 1 1705
box -2 -3 10 103
use OAI21X1  OAI21X1_133
timestamp 1696145522
transform 1 0 1004 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_270
timestamp 1696145522
transform 1 0 1036 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_246
timestamp 1696145522
transform -1 0 1092 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_320
timestamp 1696145522
transform -1 0 1116 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_302
timestamp 1696145522
transform -1 0 1148 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_128
timestamp 1696145522
transform 1 0 1148 0 1 1705
box -2 -3 26 103
use INVX1  INVX1_284
timestamp 1696145522
transform -1 0 1188 0 1 1705
box -2 -3 18 103
use NOR2X1  NOR2X1_222
timestamp 1696145522
transform -1 0 1212 0 1 1705
box -2 -3 26 103
use MUX2X1  MUX2X1_73
timestamp 1696145522
transform 1 0 1212 0 1 1705
box -2 -3 50 103
use NOR2X1  NOR2X1_316
timestamp 1696145522
transform -1 0 1284 0 1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_589
timestamp 1696145522
transform 1 0 1284 0 1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_315
timestamp 1696145522
transform -1 0 1332 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_569
timestamp 1696145522
transform 1 0 1332 0 1 1705
box -2 -3 34 103
use MUX2X1  MUX2X1_57
timestamp 1696145522
transform 1 0 1364 0 1 1705
box -2 -3 50 103
use OAI21X1  OAI21X1_735
timestamp 1696145522
transform 1 0 1412 0 1 1705
box -2 -3 34 103
use NAND3X1  NAND3X1_36
timestamp 1696145522
transform -1 0 1476 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_633
timestamp 1696145522
transform 1 0 1476 0 1 1705
box -2 -3 34 103
use FILL  FILL_17_2_0
timestamp 1696145522
transform 1 0 1508 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_2_1
timestamp 1696145522
transform 1 0 1516 0 1 1705
box -2 -3 10 103
use OAI21X1  OAI21X1_632
timestamp 1696145522
transform 1 0 1524 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_427
timestamp 1696145522
transform 1 0 1556 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_581
timestamp 1696145522
transform 1 0 1588 0 1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_229
timestamp 1696145522
transform 1 0 1620 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_494
timestamp 1696145522
transform -1 0 1676 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_903
timestamp 1696145522
transform 1 0 1676 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_580
timestamp 1696145522
transform -1 0 1740 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_917
timestamp 1696145522
transform 1 0 1740 0 1 1705
box -2 -3 34 103
use OAI22X1  OAI22X1_35
timestamp 1696145522
transform 1 0 1772 0 1 1705
box -2 -3 42 103
use NOR2X1  NOR2X1_372
timestamp 1696145522
transform 1 0 1812 0 1 1705
box -2 -3 26 103
use OAI22X1  OAI22X1_34
timestamp 1696145522
transform -1 0 1876 0 1 1705
box -2 -3 42 103
use AOI21X1  AOI21X1_221
timestamp 1696145522
transform -1 0 1908 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_911
timestamp 1696145522
transform -1 0 1940 0 1 1705
box -2 -3 34 103
use INVX1  INVX1_234
timestamp 1696145522
transform 1 0 1940 0 1 1705
box -2 -3 18 103
use BUFX4  BUFX4_169
timestamp 1696145522
transform -1 0 1988 0 1 1705
box -2 -3 34 103
use AND2X2  AND2X2_3
timestamp 1696145522
transform 1 0 1988 0 1 1705
box -2 -3 34 103
use FILL  FILL_17_3_0
timestamp 1696145522
transform 1 0 2020 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_3_1
timestamp 1696145522
transform 1 0 2028 0 1 1705
box -2 -3 10 103
use OAI22X1  OAI22X1_12
timestamp 1696145522
transform 1 0 2036 0 1 1705
box -2 -3 42 103
use AOI21X1  AOI21X1_335
timestamp 1696145522
transform 1 0 2076 0 1 1705
box -2 -3 34 103
use INVX1  INVX1_172
timestamp 1696145522
transform -1 0 2124 0 1 1705
box -2 -3 18 103
use NAND2X1  NAND2X1_464
timestamp 1696145522
transform -1 0 2148 0 1 1705
box -2 -3 26 103
use INVX1  INVX1_250
timestamp 1696145522
transform 1 0 2148 0 1 1705
box -2 -3 18 103
use OAI21X1  OAI21X1_888
timestamp 1696145522
transform 1 0 2164 0 1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_383
timestamp 1696145522
transform -1 0 2228 0 1 1705
box -2 -3 34 103
use INVX1  INVX1_133
timestamp 1696145522
transform 1 0 2228 0 1 1705
box -2 -3 18 103
use OAI21X1  OAI21X1_304
timestamp 1696145522
transform 1 0 2244 0 1 1705
box -2 -3 34 103
use OAI21X1  OAI21X1_303
timestamp 1696145522
transform 1 0 2276 0 1 1705
box -2 -3 34 103
use INVX1  INVX1_74
timestamp 1696145522
transform -1 0 2324 0 1 1705
box -2 -3 18 103
use BUFX4  BUFX4_88
timestamp 1696145522
transform -1 0 2356 0 1 1705
box -2 -3 34 103
use AND2X2  AND2X2_55
timestamp 1696145522
transform 1 0 2356 0 1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_156
timestamp 1696145522
transform -1 0 2420 0 1 1705
box -2 -3 34 103
use BUFX4  BUFX4_171
timestamp 1696145522
transform -1 0 2452 0 1 1705
box -2 -3 34 103
use INVX1  INVX1_296
timestamp 1696145522
transform 1 0 2452 0 1 1705
box -2 -3 18 103
use INVX8  INVX8_18
timestamp 1696145522
transform 1 0 2468 0 1 1705
box -2 -3 42 103
use INVX1  INVX1_176
timestamp 1696145522
transform 1 0 2508 0 1 1705
box -2 -3 18 103
use FILL  FILL_17_4_0
timestamp 1696145522
transform 1 0 2524 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_4_1
timestamp 1696145522
transform 1 0 2532 0 1 1705
box -2 -3 10 103
use AOI21X1  AOI21X1_142
timestamp 1696145522
transform 1 0 2540 0 1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_426
timestamp 1696145522
transform -1 0 2596 0 1 1705
box -2 -3 26 103
use INVX8  INVX8_10
timestamp 1696145522
transform 1 0 2596 0 1 1705
box -2 -3 42 103
use NOR2X1  NOR2X1_72
timestamp 1696145522
transform 1 0 2636 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_428
timestamp 1696145522
transform -1 0 2692 0 1 1705
box -2 -3 34 103
use NOR2X1  NOR2X1_44
timestamp 1696145522
transform 1 0 2692 0 1 1705
box -2 -3 26 103
use INVX1  INVX1_27
timestamp 1696145522
transform 1 0 2716 0 1 1705
box -2 -3 18 103
use INVX2  INVX2_37
timestamp 1696145522
transform 1 0 2732 0 1 1705
box -2 -3 18 103
use INVX1  INVX1_35
timestamp 1696145522
transform 1 0 2748 0 1 1705
box -2 -3 18 103
use NOR2X1  NOR2X1_78
timestamp 1696145522
transform -1 0 2788 0 1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_45
timestamp 1696145522
transform -1 0 2812 0 1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_85
timestamp 1696145522
transform -1 0 2836 0 1 1705
box -2 -3 26 103
use INVX2  INVX2_33
timestamp 1696145522
transform -1 0 2852 0 1 1705
box -2 -3 18 103
use NOR2X1  NOR2X1_43
timestamp 1696145522
transform 1 0 2852 0 1 1705
box -2 -3 26 103
use NAND2X1  NAND2X1_639
timestamp 1696145522
transform 1 0 2876 0 1 1705
box -2 -3 26 103
use AOI22X1  AOI22X1_52
timestamp 1696145522
transform -1 0 2940 0 1 1705
box -2 -3 42 103
use NOR2X1  NOR2X1_12
timestamp 1696145522
transform 1 0 2940 0 1 1705
box -2 -3 26 103
use OR2X2  OR2X2_49
timestamp 1696145522
transform 1 0 2964 0 1 1705
box -2 -3 34 103
use XOR2X1  XOR2X1_1
timestamp 1696145522
transform 1 0 2996 0 1 1705
box -2 -3 58 103
use FILL  FILL_17_5_0
timestamp 1696145522
transform -1 0 3060 0 1 1705
box -2 -3 10 103
use FILL  FILL_17_5_1
timestamp 1696145522
transform -1 0 3068 0 1 1705
box -2 -3 10 103
use NOR2X1  NOR2X1_53
timestamp 1696145522
transform -1 0 3092 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_1
timestamp 1696145522
transform -1 0 3124 0 1 1705
box -2 -3 34 103
use INVX1  INVX1_3
timestamp 1696145522
transform 1 0 3124 0 1 1705
box -2 -3 18 103
use OAI21X1  OAI21X1_646
timestamp 1696145522
transform 1 0 3140 0 1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_21
timestamp 1696145522
transform 1 0 3172 0 1 1705
box -2 -3 34 103
use NAND2X1  NAND2X1_4
timestamp 1696145522
transform -1 0 3228 0 1 1705
box -2 -3 26 103
use INVX1  INVX1_9
timestamp 1696145522
transform -1 0 3244 0 1 1705
box -2 -3 18 103
use NOR2X1  NOR2X1_4
timestamp 1696145522
transform 1 0 3244 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_906
timestamp 1696145522
transform 1 0 3268 0 1 1705
box -2 -3 34 103
use XNOR2X1  XNOR2X1_10
timestamp 1696145522
transform 1 0 3300 0 1 1705
box -2 -3 58 103
use NAND2X1  NAND2X1_60
timestamp 1696145522
transform -1 0 3380 0 1 1705
box -2 -3 26 103
use OAI21X1  OAI21X1_904
timestamp 1696145522
transform -1 0 3412 0 1 1705
box -2 -3 34 103
use CLKBUF1  CLKBUF1_6
timestamp 1696145522
transform 1 0 3412 0 1 1705
box -2 -3 74 103
use OAI21X1  OAI21X1_636
timestamp 1696145522
transform 1 0 3484 0 1 1705
box -2 -3 34 103
use AOI21X1  AOI21X1_387
timestamp 1696145522
transform -1 0 3548 0 1 1705
box -2 -3 34 103
use INVX1  INVX1_330
timestamp 1696145522
transform -1 0 3564 0 1 1705
box -2 -3 18 103
use BUFX4  BUFX4_70
timestamp 1696145522
transform -1 0 36 0 -1 1905
box -2 -3 34 103
use MUX2X1  MUX2X1_62
timestamp 1696145522
transform -1 0 84 0 -1 1905
box -2 -3 50 103
use INVX1  INVX1_227
timestamp 1696145522
transform -1 0 100 0 -1 1905
box -2 -3 18 103
use OAI21X1  OAI21X1_197
timestamp 1696145522
transform -1 0 132 0 -1 1905
box -2 -3 34 103
use INVX1  INVX1_95
timestamp 1696145522
transform -1 0 148 0 -1 1905
box -2 -3 18 103
use NAND2X1  NAND2X1_455
timestamp 1696145522
transform 1 0 148 0 -1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_513
timestamp 1696145522
transform -1 0 204 0 -1 1905
box -2 -3 34 103
use INVX1  INVX1_213
timestamp 1696145522
transform -1 0 220 0 -1 1905
box -2 -3 18 103
use MUX2X1  MUX2X1_61
timestamp 1696145522
transform 1 0 220 0 -1 1905
box -2 -3 50 103
use OAI21X1  OAI21X1_527
timestamp 1696145522
transform -1 0 300 0 -1 1905
box -2 -3 34 103
use MUX2X1  MUX2X1_41
timestamp 1696145522
transform 1 0 300 0 -1 1905
box -2 -3 50 103
use NAND2X1  NAND2X1_472
timestamp 1696145522
transform 1 0 348 0 -1 1905
box -2 -3 26 103
use MUX2X1  MUX2X1_45
timestamp 1696145522
transform 1 0 372 0 -1 1905
box -2 -3 50 103
use MUX2X1  MUX2X1_51
timestamp 1696145522
transform -1 0 468 0 -1 1905
box -2 -3 50 103
use INVX1  INVX1_121
timestamp 1696145522
transform -1 0 484 0 -1 1905
box -2 -3 18 103
use FILL  FILL_18_0_0
timestamp 1696145522
transform -1 0 492 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_0_1
timestamp 1696145522
transform -1 0 500 0 -1 1905
box -2 -3 10 103
use INVX1  INVX1_206
timestamp 1696145522
transform -1 0 516 0 -1 1905
box -2 -3 18 103
use INVX1  INVX1_174
timestamp 1696145522
transform -1 0 532 0 -1 1905
box -2 -3 18 103
use OAI21X1  OAI21X1_441
timestamp 1696145522
transform 1 0 532 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_229
timestamp 1696145522
transform -1 0 596 0 -1 1905
box -2 -3 34 103
use INVX1  INVX1_165
timestamp 1696145522
transform -1 0 612 0 -1 1905
box -2 -3 18 103
use NAND2X1  NAND2X1_250
timestamp 1696145522
transform 1 0 612 0 -1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_219
timestamp 1696145522
transform -1 0 668 0 -1 1905
box -2 -3 34 103
use INVX1  INVX1_61
timestamp 1696145522
transform -1 0 684 0 -1 1905
box -2 -3 18 103
use OAI21X1  OAI21X1_177
timestamp 1696145522
transform -1 0 716 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_319
timestamp 1696145522
transform -1 0 740 0 -1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_210
timestamp 1696145522
transform 1 0 740 0 -1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_124
timestamp 1696145522
transform 1 0 764 0 -1 1905
box -2 -3 26 103
use MUX2X1  MUX2X1_30
timestamp 1696145522
transform 1 0 788 0 -1 1905
box -2 -3 50 103
use OAI21X1  OAI21X1_245
timestamp 1696145522
transform 1 0 836 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_269
timestamp 1696145522
transform 1 0 868 0 -1 1905
box -2 -3 26 103
use INVX1  INVX1_50
timestamp 1696145522
transform -1 0 908 0 -1 1905
box -2 -3 18 103
use OAI21X1  OAI21X1_84
timestamp 1696145522
transform 1 0 908 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_135
timestamp 1696145522
transform 1 0 940 0 -1 1905
box -2 -3 26 103
use INVX1  INVX1_69
timestamp 1696145522
transform 1 0 964 0 -1 1905
box -2 -3 18 103
use NAND2X1  NAND2X1_177
timestamp 1696145522
transform -1 0 1004 0 -1 1905
box -2 -3 26 103
use FILL  FILL_18_1_0
timestamp 1696145522
transform 1 0 1004 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_1_1
timestamp 1696145522
transform 1 0 1012 0 -1 1905
box -2 -3 10 103
use OAI21X1  OAI21X1_300
timestamp 1696145522
transform 1 0 1020 0 -1 1905
box -2 -3 34 103
use INVX1  INVX1_70
timestamp 1696145522
transform -1 0 1068 0 -1 1905
box -2 -3 18 103
use NAND2X1  NAND2X1_292
timestamp 1696145522
transform -1 0 1092 0 -1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_266
timestamp 1696145522
transform -1 0 1124 0 -1 1905
box -2 -3 34 103
use MUX2X1  MUX2X1_24
timestamp 1696145522
transform 1 0 1124 0 -1 1905
box -2 -3 50 103
use MUX2X1  MUX2X1_103
timestamp 1696145522
transform 1 0 1172 0 -1 1905
box -2 -3 50 103
use MUX2X1  MUX2X1_71
timestamp 1696145522
transform -1 0 1268 0 -1 1905
box -2 -3 50 103
use MUX2X1  MUX2X1_20
timestamp 1696145522
transform 1 0 1268 0 -1 1905
box -2 -3 50 103
use NAND2X1  NAND2X1_92
timestamp 1696145522
transform 1 0 1316 0 -1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_485
timestamp 1696145522
transform -1 0 1364 0 -1 1905
box -2 -3 26 103
use AOI21X1  AOI21X1_254
timestamp 1696145522
transform 1 0 1364 0 -1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_255
timestamp 1696145522
transform 1 0 1396 0 -1 1905
box -2 -3 34 103
use MUX2X1  MUX2X1_79
timestamp 1696145522
transform 1 0 1428 0 -1 1905
box -2 -3 50 103
use AOI21X1  AOI21X1_256
timestamp 1696145522
transform -1 0 1508 0 -1 1905
box -2 -3 34 103
use FILL  FILL_18_2_0
timestamp 1696145522
transform 1 0 1508 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_2_1
timestamp 1696145522
transform 1 0 1516 0 -1 1905
box -2 -3 10 103
use AOI21X1  AOI21X1_236
timestamp 1696145522
transform 1 0 1524 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_588
timestamp 1696145522
transform 1 0 1556 0 -1 1905
box -2 -3 34 103
use AND2X2  AND2X2_75
timestamp 1696145522
transform 1 0 1588 0 -1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_237
timestamp 1696145522
transform 1 0 1620 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_515
timestamp 1696145522
transform -1 0 1676 0 -1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_939
timestamp 1696145522
transform 1 0 1676 0 -1 1905
box -2 -3 34 103
use OAI22X1  OAI22X1_38
timestamp 1696145522
transform -1 0 1748 0 -1 1905
box -2 -3 42 103
use NAND2X1  NAND2X1_496
timestamp 1696145522
transform -1 0 1772 0 -1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_505
timestamp 1696145522
transform 1 0 1772 0 -1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_926
timestamp 1696145522
transform 1 0 1796 0 -1 1905
box -2 -3 34 103
use OAI22X1  OAI22X1_36
timestamp 1696145522
transform -1 0 1868 0 -1 1905
box -2 -3 42 103
use NAND2X1  NAND2X1_374
timestamp 1696145522
transform -1 0 1892 0 -1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_503
timestamp 1696145522
transform 1 0 1892 0 -1 1905
box -2 -3 26 103
use AOI21X1  AOI21X1_234
timestamp 1696145522
transform 1 0 1916 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_946
timestamp 1696145522
transform 1 0 1948 0 -1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_260
timestamp 1696145522
transform -1 0 2012 0 -1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_509
timestamp 1696145522
transform -1 0 2036 0 -1 1905
box -2 -3 26 103
use FILL  FILL_18_3_0
timestamp 1696145522
transform -1 0 2044 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_3_1
timestamp 1696145522
transform -1 0 2052 0 -1 1905
box -2 -3 10 103
use AOI21X1  AOI21X1_129
timestamp 1696145522
transform -1 0 2084 0 -1 1905
box -2 -3 34 103
use BUFX4  BUFX4_174
timestamp 1696145522
transform -1 0 2116 0 -1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_253
timestamp 1696145522
transform -1 0 2148 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_603
timestamp 1696145522
transform 1 0 2148 0 -1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_194
timestamp 1696145522
transform -1 0 2212 0 -1 1905
box -2 -3 34 103
use OR2X2  OR2X2_14
timestamp 1696145522
transform -1 0 2244 0 -1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_88
timestamp 1696145522
transform -1 0 2276 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_315
timestamp 1696145522
transform -1 0 2300 0 -1 1905
box -2 -3 26 103
use AOI21X1  AOI21X1_42
timestamp 1696145522
transform 1 0 2300 0 -1 1905
box -2 -3 34 103
use INVX4  INVX4_20
timestamp 1696145522
transform 1 0 2332 0 -1 1905
box -2 -3 26 103
use BUFX4  BUFX4_8
timestamp 1696145522
transform -1 0 2388 0 -1 1905
box -2 -3 34 103
use INVX8  INVX8_12
timestamp 1696145522
transform 1 0 2388 0 -1 1905
box -2 -3 42 103
use INVX2  INVX2_8
timestamp 1696145522
transform 1 0 2428 0 -1 1905
box -2 -3 18 103
use INVX8  INVX8_7
timestamp 1696145522
transform 1 0 2444 0 -1 1905
box -2 -3 42 103
use INVX4  INVX4_18
timestamp 1696145522
transform 1 0 2484 0 -1 1905
box -2 -3 26 103
use OR2X2  OR2X2_23
timestamp 1696145522
transform -1 0 2540 0 -1 1905
box -2 -3 34 103
use FILL  FILL_18_4_0
timestamp 1696145522
transform -1 0 2548 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_4_1
timestamp 1696145522
transform -1 0 2556 0 -1 1905
box -2 -3 10 103
use NAND3X1  NAND3X1_22
timestamp 1696145522
transform -1 0 2588 0 -1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_10
timestamp 1696145522
transform 1 0 2588 0 -1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_74
timestamp 1696145522
transform 1 0 2620 0 -1 1905
box -2 -3 26 103
use INVX2  INVX2_34
timestamp 1696145522
transform 1 0 2644 0 -1 1905
box -2 -3 18 103
use NOR2X1  NOR2X1_71
timestamp 1696145522
transform 1 0 2660 0 -1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_413
timestamp 1696145522
transform 1 0 2684 0 -1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_675
timestamp 1696145522
transform 1 0 2708 0 -1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_296
timestamp 1696145522
transform 1 0 2740 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_556
timestamp 1696145522
transform -1 0 2796 0 -1 1905
box -2 -3 26 103
use INVX2  INVX2_36
timestamp 1696145522
transform -1 0 2812 0 -1 1905
box -2 -3 18 103
use NOR2X1  NOR2X1_73
timestamp 1696145522
transform 1 0 2812 0 -1 1905
box -2 -3 26 103
use AOI21X1  AOI21X1_50
timestamp 1696145522
transform 1 0 2836 0 -1 1905
box -2 -3 34 103
use INVX1  INVX1_43
timestamp 1696145522
transform -1 0 2884 0 -1 1905
box -2 -3 18 103
use AND2X2  AND2X2_1
timestamp 1696145522
transform -1 0 2916 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_191
timestamp 1696145522
transform -1 0 2940 0 -1 1905
box -2 -3 26 103
use XNOR2X1  XNOR2X1_46
timestamp 1696145522
transform 1 0 2940 0 -1 1905
box -2 -3 58 103
use AOI21X1  AOI21X1_281
timestamp 1696145522
transform 1 0 2996 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_205
timestamp 1696145522
transform -1 0 3052 0 -1 1905
box -2 -3 26 103
use FILL  FILL_18_5_0
timestamp 1696145522
transform 1 0 3052 0 -1 1905
box -2 -3 10 103
use FILL  FILL_18_5_1
timestamp 1696145522
transform 1 0 3060 0 -1 1905
box -2 -3 10 103
use AOI21X1  AOI21X1_32
timestamp 1696145522
transform 1 0 3068 0 -1 1905
box -2 -3 34 103
use INVX1  INVX1_31
timestamp 1696145522
transform -1 0 3116 0 -1 1905
box -2 -3 18 103
use OAI21X1  OAI21X1_651
timestamp 1696145522
transform -1 0 3148 0 -1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_65
timestamp 1696145522
transform 1 0 3148 0 -1 1905
box -2 -3 26 103
use XNOR2X1  XNOR2X1_11
timestamp 1696145522
transform 1 0 3172 0 -1 1905
box -2 -3 58 103
use AOI21X1  AOI21X1_390
timestamp 1696145522
transform -1 0 3260 0 -1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_907
timestamp 1696145522
transform -1 0 3292 0 -1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_25
timestamp 1696145522
transform 1 0 3292 0 -1 1905
box -2 -3 98 103
use OAI21X1  OAI21X1_905
timestamp 1696145522
transform 1 0 3388 0 -1 1905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_23
timestamp 1696145522
transform 1 0 3420 0 -1 1905
box -2 -3 98 103
use INVX1  INVX1_277
timestamp 1696145522
transform -1 0 3532 0 -1 1905
box -2 -3 18 103
use BUFX2  BUFX2_25
timestamp 1696145522
transform 1 0 3532 0 -1 1905
box -2 -3 26 103
use FILL  FILL_19_1
timestamp 1696145522
transform -1 0 3564 0 -1 1905
box -2 -3 10 103
use OAI21X1  OAI21X1_614
timestamp 1696145522
transform 1 0 4 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_518
timestamp 1696145522
transform 1 0 36 0 1 1905
box -2 -3 26 103
use INVX1  INVX1_254
timestamp 1696145522
transform -1 0 76 0 1 1905
box -2 -3 18 103
use OAI21X1  OAI21X1_232
timestamp 1696145522
transform -1 0 108 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_168
timestamp 1696145522
transform -1 0 132 0 1 1905
box -2 -3 26 103
use MUX2X1  MUX2X1_60
timestamp 1696145522
transform -1 0 180 0 1 1905
box -2 -3 50 103
use OAI21X1  OAI21X1_628
timestamp 1696145522
transform 1 0 180 0 1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_274
timestamp 1696145522
transform -1 0 244 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_230
timestamp 1696145522
transform -1 0 268 0 1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_440
timestamp 1696145522
transform 1 0 268 0 1 1905
box -2 -3 26 103
use INVX1  INVX1_217
timestamp 1696145522
transform -1 0 308 0 1 1905
box -2 -3 18 103
use MUX2X1  MUX2X1_66
timestamp 1696145522
transform -1 0 356 0 1 1905
box -2 -3 50 103
use NAND2X1  NAND2X1_467
timestamp 1696145522
transform 1 0 356 0 1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_504
timestamp 1696145522
transform -1 0 404 0 1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_493
timestamp 1696145522
transform 1 0 404 0 1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_171
timestamp 1696145522
transform -1 0 452 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_127
timestamp 1696145522
transform -1 0 484 0 1 1905
box -2 -3 34 103
use FILL  FILL_19_0_0
timestamp 1696145522
transform -1 0 492 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_0_1
timestamp 1696145522
transform -1 0 500 0 1 1905
box -2 -3 10 103
use OAI21X1  OAI21X1_468
timestamp 1696145522
transform -1 0 532 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_65
timestamp 1696145522
transform -1 0 564 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_258
timestamp 1696145522
transform -1 0 588 0 1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_414
timestamp 1696145522
transform -1 0 612 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_323
timestamp 1696145522
transform -1 0 644 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_349
timestamp 1696145522
transform 1 0 644 0 1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_82
timestamp 1696145522
transform -1 0 700 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_175
timestamp 1696145522
transform 1 0 700 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_176
timestamp 1696145522
transform -1 0 756 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_107
timestamp 1696145522
transform 1 0 756 0 1 1905
box -2 -3 34 103
use BUFX4  BUFX4_68
timestamp 1696145522
transform 1 0 788 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_132
timestamp 1696145522
transform -1 0 852 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_230
timestamp 1696145522
transform 1 0 852 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_132
timestamp 1696145522
transform -1 0 908 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_81
timestamp 1696145522
transform -1 0 940 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_217
timestamp 1696145522
transform 1 0 940 0 1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_216
timestamp 1696145522
transform -1 0 988 0 1 1905
box -2 -3 26 103
use FILL  FILL_19_1_0
timestamp 1696145522
transform -1 0 996 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_1_1
timestamp 1696145522
transform -1 0 1004 0 1 1905
box -2 -3 10 103
use OAI21X1  OAI21X1_183
timestamp 1696145522
transform -1 0 1036 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_317
timestamp 1696145522
transform -1 0 1060 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_136
timestamp 1696145522
transform -1 0 1092 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_226
timestamp 1696145522
transform 1 0 1092 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_255
timestamp 1696145522
transform -1 0 1148 0 1 1905
box -2 -3 26 103
use NAND2X1  NAND2X1_581
timestamp 1696145522
transform 1 0 1148 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_722
timestamp 1696145522
transform -1 0 1204 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_141
timestamp 1696145522
transform 1 0 1204 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_184
timestamp 1696145522
transform -1 0 1260 0 1 1905
box -2 -3 26 103
use OAI21X1  OAI21X1_677
timestamp 1696145522
transform 1 0 1260 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_43
timestamp 1696145522
transform 1 0 1292 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_733
timestamp 1696145522
transform 1 0 1324 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_551
timestamp 1696145522
transform -1 0 1388 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_607
timestamp 1696145522
transform -1 0 1420 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_590
timestamp 1696145522
transform 1 0 1420 0 1 1905
box -2 -3 26 103
use AOI21X1  AOI21X1_213
timestamp 1696145522
transform -1 0 1476 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_606
timestamp 1696145522
transform -1 0 1508 0 1 1905
box -2 -3 34 103
use FILL  FILL_19_2_0
timestamp 1696145522
transform -1 0 1516 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_2_1
timestamp 1696145522
transform -1 0 1524 0 1 1905
box -2 -3 10 103
use OAI21X1  OAI21X1_550
timestamp 1696145522
transform -1 0 1556 0 1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_206
timestamp 1696145522
transform -1 0 1588 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_595
timestamp 1696145522
transform 1 0 1588 0 1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_244
timestamp 1696145522
transform -1 0 1652 0 1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_222
timestamp 1696145522
transform 1 0 1652 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_587
timestamp 1696145522
transform -1 0 1716 0 1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_34
timestamp 1696145522
transform 1 0 1716 0 1 1905
box -2 -3 34 103
use OR2X2  OR2X2_32
timestamp 1696145522
transform -1 0 1780 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_618
timestamp 1696145522
transform -1 0 1812 0 1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_261
timestamp 1696145522
transform -1 0 1844 0 1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_17
timestamp 1696145522
transform 1 0 1844 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_487
timestamp 1696145522
transform -1 0 1908 0 1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_169
timestamp 1696145522
transform -1 0 1940 0 1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_19
timestamp 1696145522
transform 1 0 1940 0 1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_98
timestamp 1696145522
transform 1 0 1972 0 1 1905
box -2 -3 26 103
use INVX1  INVX1_72
timestamp 1696145522
transform 1 0 1996 0 1 1905
box -2 -3 18 103
use FILL  FILL_19_3_0
timestamp 1696145522
transform 1 0 2012 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_3_1
timestamp 1696145522
transform 1 0 2020 0 1 1905
box -2 -3 10 103
use OAI21X1  OAI21X1_146
timestamp 1696145522
transform 1 0 2028 0 1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_161
timestamp 1696145522
transform 1 0 2060 0 1 1905
box -2 -3 26 103
use NOR2X1  NOR2X1_175
timestamp 1696145522
transform -1 0 2108 0 1 1905
box -2 -3 26 103
use OR2X2  OR2X2_19
timestamp 1696145522
transform -1 0 2140 0 1 1905
box -2 -3 34 103
use INVX1  INVX1_145
timestamp 1696145522
transform 1 0 2140 0 1 1905
box -2 -3 18 103
use OAI21X1  OAI21X1_367
timestamp 1696145522
transform 1 0 2156 0 1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_13
timestamp 1696145522
transform 1 0 2188 0 1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_87
timestamp 1696145522
transform -1 0 2252 0 1 1905
box -2 -3 34 103
use NAND3X1  NAND3X1_12
timestamp 1696145522
transform -1 0 2284 0 1 1905
box -2 -3 34 103
use OR2X2  OR2X2_26
timestamp 1696145522
transform 1 0 2284 0 1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_167
timestamp 1696145522
transform -1 0 2340 0 1 1905
box -2 -3 26 103
use AND2X2  AND2X2_8
timestamp 1696145522
transform 1 0 2340 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_148
timestamp 1696145522
transform 1 0 2372 0 1 1905
box -2 -3 34 103
use BUFX4  BUFX4_59
timestamp 1696145522
transform 1 0 2404 0 1 1905
box -2 -3 34 103
use BUFX4  BUFX4_62
timestamp 1696145522
transform -1 0 2468 0 1 1905
box -2 -3 34 103
use INVX2  INVX2_32
timestamp 1696145522
transform -1 0 2484 0 1 1905
box -2 -3 18 103
use NOR2X1  NOR2X1_224
timestamp 1696145522
transform -1 0 2508 0 1 1905
box -2 -3 26 103
use BUFX4  BUFX4_27
timestamp 1696145522
transform -1 0 2540 0 1 1905
box -2 -3 34 103
use FILL  FILL_19_4_0
timestamp 1696145522
transform 1 0 2540 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_4_1
timestamp 1696145522
transform 1 0 2548 0 1 1905
box -2 -3 10 103
use OAI21X1  OAI21X1_950
timestamp 1696145522
transform 1 0 2556 0 1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_148
timestamp 1696145522
transform 1 0 2588 0 1 1905
box -2 -3 26 103
use BUFX4  BUFX4_148
timestamp 1696145522
transform 1 0 2612 0 1 1905
box -2 -3 34 103
use BUFX4  BUFX4_106
timestamp 1696145522
transform 1 0 2644 0 1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_295
timestamp 1696145522
transform 1 0 2676 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_538
timestamp 1696145522
transform -1 0 2732 0 1 1905
box -2 -3 26 103
use NAND3X1  NAND3X1_72
timestamp 1696145522
transform -1 0 2764 0 1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_397
timestamp 1696145522
transform 1 0 2764 0 1 1905
box -2 -3 34 103
use INVX1  INVX1_323
timestamp 1696145522
transform 1 0 2796 0 1 1905
box -2 -3 18 103
use AOI21X1  AOI21X1_393
timestamp 1696145522
transform 1 0 2812 0 1 1905
box -2 -3 34 103
use NAND2X1  NAND2X1_198
timestamp 1696145522
transform 1 0 2844 0 1 1905
box -2 -3 26 103
use AOI21X1  AOI21X1_15
timestamp 1696145522
transform 1 0 2868 0 1 1905
box -2 -3 34 103
use INVX1  INVX1_10
timestamp 1696145522
transform -1 0 2916 0 1 1905
box -2 -3 18 103
use AOI21X1  AOI21X1_61
timestamp 1696145522
transform 1 0 2916 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_655
timestamp 1696145522
transform -1 0 2980 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_168
timestamp 1696145522
transform 1 0 2980 0 1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_499
timestamp 1696145522
transform -1 0 3036 0 1 1905
box -2 -3 26 103
use FILL  FILL_19_5_0
timestamp 1696145522
transform 1 0 3036 0 1 1905
box -2 -3 10 103
use FILL  FILL_19_5_1
timestamp 1696145522
transform 1 0 3044 0 1 1905
box -2 -3 10 103
use BUFX4  BUFX4_31
timestamp 1696145522
transform 1 0 3052 0 1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_57
timestamp 1696145522
transform 1 0 3084 0 1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_122
timestamp 1696145522
transform 1 0 3116 0 1 1905
box -2 -3 26 103
use AOI21X1  AOI21X1_394
timestamp 1696145522
transform 1 0 3140 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_909
timestamp 1696145522
transform 1 0 3172 0 1 1905
box -2 -3 34 103
use AOI21X1  AOI21X1_398
timestamp 1696145522
transform 1 0 3204 0 1 1905
box -2 -3 34 103
use OAI21X1  OAI21X1_174
timestamp 1696145522
transform 1 0 3236 0 1 1905
box -2 -3 34 103
use AOI22X1  AOI22X1_54
timestamp 1696145522
transform -1 0 3308 0 1 1905
box -2 -3 42 103
use NOR2X1  NOR2X1_498
timestamp 1696145522
transform 1 0 3308 0 1 1905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_24
timestamp 1696145522
transform 1 0 3332 0 1 1905
box -2 -3 98 103
use INVX1  INVX1_276
timestamp 1696145522
transform 1 0 3428 0 1 1905
box -2 -3 18 103
use NAND3X1  NAND3X1_51
timestamp 1696145522
transform 1 0 3444 0 1 1905
box -2 -3 34 103
use NOR2X1  NOR2X1_405
timestamp 1696145522
transform -1 0 3500 0 1 1905
box -2 -3 26 103
use BUFX2  BUFX2_26
timestamp 1696145522
transform 1 0 3500 0 1 1905
box -2 -3 26 103
use BUFX2  BUFX2_27
timestamp 1696145522
transform 1 0 3524 0 1 1905
box -2 -3 26 103
use FILL  FILL_20_1
timestamp 1696145522
transform 1 0 3548 0 1 1905
box -2 -3 10 103
use FILL  FILL_20_2
timestamp 1696145522
transform 1 0 3556 0 1 1905
box -2 -3 10 103
use NAND2X1  NAND2X1_509
timestamp 1696145522
transform 1 0 4 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_592
timestamp 1696145522
transform -1 0 60 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_262
timestamp 1696145522
transform 1 0 60 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_613
timestamp 1696145522
transform 1 0 84 0 -1 2105
box -2 -3 34 103
use INVX1  INVX1_131
timestamp 1696145522
transform -1 0 132 0 -1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_557
timestamp 1696145522
transform -1 0 164 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_124
timestamp 1696145522
transform 1 0 164 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_48
timestamp 1696145522
transform -1 0 228 0 -1 2105
box -2 -3 34 103
use INVX1  INVX1_41
timestamp 1696145522
transform -1 0 244 0 -1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_512
timestamp 1696145522
transform -1 0 276 0 -1 2105
box -2 -3 34 103
use INVX1  INVX1_115
timestamp 1696145522
transform -1 0 292 0 -1 2105
box -2 -3 18 103
use INVX1  INVX1_178
timestamp 1696145522
transform -1 0 308 0 -1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_199
timestamp 1696145522
transform 1 0 308 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_535
timestamp 1696145522
transform 1 0 340 0 -1 2105
box -2 -3 34 103
use MUX2X1  MUX2X1_22
timestamp 1696145522
transform 1 0 372 0 -1 2105
box -2 -3 50 103
use NAND2X1  NAND2X1_116
timestamp 1696145522
transform -1 0 444 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_62
timestamp 1696145522
transform 1 0 444 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_111
timestamp 1696145522
transform -1 0 500 0 -1 2105
box -2 -3 26 103
use FILL  FILL_20_0_0
timestamp 1696145522
transform 1 0 500 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_0_1
timestamp 1696145522
transform 1 0 508 0 -1 2105
box -2 -3 10 103
use OAI21X1  OAI21X1_492
timestamp 1696145522
transform 1 0 516 0 -1 2105
box -2 -3 34 103
use INVX1  INVX1_47
timestamp 1696145522
transform -1 0 564 0 -1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_413
timestamp 1696145522
transform -1 0 596 0 -1 2105
box -2 -3 34 103
use MUX2X1  MUX2X1_23
timestamp 1696145522
transform 1 0 596 0 -1 2105
box -2 -3 50 103
use NAND2X1  NAND2X1_336
timestamp 1696145522
transform 1 0 644 0 -1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_298
timestamp 1696145522
transform 1 0 668 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_276
timestamp 1696145522
transform -1 0 724 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_218
timestamp 1696145522
transform 1 0 724 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_176
timestamp 1696145522
transform 1 0 756 0 -1 2105
box -2 -3 34 103
use INVX1  INVX1_49
timestamp 1696145522
transform 1 0 788 0 -1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_72
timestamp 1696145522
transform 1 0 804 0 -1 2105
box -2 -3 34 103
use INVX1  INVX1_87
timestamp 1696145522
transform 1 0 836 0 -1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_182
timestamp 1696145522
transform 1 0 852 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_215
timestamp 1696145522
transform -1 0 908 0 -1 2105
box -2 -3 26 103
use INVX1  INVX1_63
timestamp 1696145522
transform -1 0 924 0 -1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_130
timestamp 1696145522
transform -1 0 956 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_224
timestamp 1696145522
transform -1 0 988 0 -1 2105
box -2 -3 34 103
use FILL  FILL_20_1_0
timestamp 1696145522
transform 1 0 988 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_1_1
timestamp 1696145522
transform 1 0 996 0 -1 2105
box -2 -3 10 103
use OAI21X1  OAI21X1_138
timestamp 1696145522
transform 1 0 1004 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_83
timestamp 1696145522
transform 1 0 1036 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_134
timestamp 1696145522
transform -1 0 1092 0 -1 2105
box -2 -3 26 103
use INVX1  INVX1_180
timestamp 1696145522
transform -1 0 1108 0 -1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_180
timestamp 1696145522
transform 1 0 1108 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_213
timestamp 1696145522
transform 1 0 1140 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_76
timestamp 1696145522
transform 1 0 1164 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_227
timestamp 1696145522
transform -1 0 1228 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_78
timestamp 1696145522
transform -1 0 1260 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_557
timestamp 1696145522
transform 1 0 1260 0 -1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_584
timestamp 1696145522
transform 1 0 1284 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_725
timestamp 1696145522
transform -1 0 1340 0 -1 2105
box -2 -3 34 103
use INVX1  INVX1_71
timestamp 1696145522
transform 1 0 1340 0 -1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_144
timestamp 1696145522
transform 1 0 1356 0 -1 2105
box -2 -3 34 103
use MUX2X1  MUX2X1_69
timestamp 1696145522
transform 1 0 1388 0 -1 2105
box -2 -3 50 103
use INVX1  INVX1_294
timestamp 1696145522
transform -1 0 1452 0 -1 2105
box -2 -3 18 103
use OAI21X1  OAI21X1_705
timestamp 1696145522
transform 1 0 1452 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_570
timestamp 1696145522
transform 1 0 1484 0 -1 2105
box -2 -3 26 103
use FILL  FILL_20_2_0
timestamp 1696145522
transform 1 0 1508 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_2_1
timestamp 1696145522
transform 1 0 1516 0 -1 2105
box -2 -3 10 103
use MUX2X1  MUX2X1_70
timestamp 1696145522
transform 1 0 1524 0 -1 2105
box -2 -3 50 103
use NAND2X1  NAND2X1_93
timestamp 1696145522
transform -1 0 1596 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_44
timestamp 1696145522
transform -1 0 1628 0 -1 2105
box -2 -3 34 103
use OR2X2  OR2X2_35
timestamp 1696145522
transform 1 0 1628 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_147
timestamp 1696145522
transform 1 0 1660 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_102
timestamp 1696145522
transform -1 0 1716 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_704
timestamp 1696145522
transform 1 0 1716 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_103
timestamp 1696145522
transform -1 0 1780 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_459
timestamp 1696145522
transform -1 0 1804 0 -1 2105
box -2 -3 26 103
use AOI21X1  AOI21X1_188
timestamp 1696145522
transform -1 0 1836 0 -1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_254
timestamp 1696145522
transform -1 0 1860 0 -1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_524
timestamp 1696145522
transform -1 0 1884 0 -1 2105
box -2 -3 26 103
use NAND3X1  NAND3X1_28
timestamp 1696145522
transform 1 0 1884 0 -1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_270
timestamp 1696145522
transform -1 0 1948 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_527
timestamp 1696145522
transform 1 0 1948 0 -1 2105
box -2 -3 26 103
use OR2X2  OR2X2_20
timestamp 1696145522
transform 1 0 1972 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_409
timestamp 1696145522
transform -1 0 2028 0 -1 2105
box -2 -3 26 103
use FILL  FILL_20_3_0
timestamp 1696145522
transform 1 0 2028 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_3_1
timestamp 1696145522
transform 1 0 2036 0 -1 2105
box -2 -3 10 103
use INVX1  INVX1_182
timestamp 1696145522
transform 1 0 2044 0 -1 2105
box -2 -3 18 103
use OR2X2  OR2X2_18
timestamp 1696145522
transform 1 0 2060 0 -1 2105
box -2 -3 34 103
use AOI22X1  AOI22X1_14
timestamp 1696145522
transform 1 0 2092 0 -1 2105
box -2 -3 42 103
use NAND3X1  NAND3X1_23
timestamp 1696145522
transform 1 0 2132 0 -1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_186
timestamp 1696145522
transform 1 0 2164 0 -1 2105
box -2 -3 26 103
use NOR2X1  NOR2X1_171
timestamp 1696145522
transform -1 0 2212 0 -1 2105
box -2 -3 26 103
use INVX2  INVX2_30
timestamp 1696145522
transform -1 0 2228 0 -1 2105
box -2 -3 18 103
use INVX8  INVX8_17
timestamp 1696145522
transform 1 0 2228 0 -1 2105
box -2 -3 42 103
use NOR2X1  NOR2X1_162
timestamp 1696145522
transform -1 0 2292 0 -1 2105
box -2 -3 26 103
use OAI22X1  OAI22X1_4
timestamp 1696145522
transform -1 0 2332 0 -1 2105
box -2 -3 42 103
use XNOR2X1  XNOR2X1_34
timestamp 1696145522
transform -1 0 2388 0 -1 2105
box -2 -3 58 103
use AOI21X1  AOI21X1_150
timestamp 1696145522
transform 1 0 2388 0 -1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_147
timestamp 1696145522
transform 1 0 2420 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_437
timestamp 1696145522
transform 1 0 2452 0 -1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_151
timestamp 1696145522
transform 1 0 2484 0 -1 2105
box -2 -3 34 103
use OR2X2  OR2X2_4
timestamp 1696145522
transform -1 0 2548 0 -1 2105
box -2 -3 34 103
use FILL  FILL_20_4_0
timestamp 1696145522
transform 1 0 2548 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_4_1
timestamp 1696145522
transform 1 0 2556 0 -1 2105
box -2 -3 10 103
use OR2X2  OR2X2_8
timestamp 1696145522
transform 1 0 2564 0 -1 2105
box -2 -3 34 103
use INVX4  INVX4_8
timestamp 1696145522
transform -1 0 2620 0 -1 2105
box -2 -3 26 103
use BUFX4  BUFX4_107
timestamp 1696145522
transform -1 0 2652 0 -1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_644
timestamp 1696145522
transform -1 0 2676 0 -1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_53
timestamp 1696145522
transform 1 0 2676 0 -1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_55
timestamp 1696145522
transform 1 0 2700 0 -1 2105
box -2 -3 26 103
use INVX1  INVX1_23
timestamp 1696145522
transform -1 0 2740 0 -1 2105
box -2 -3 18 103
use NAND2X1  NAND2X1_54
timestamp 1696145522
transform -1 0 2764 0 -1 2105
box -2 -3 26 103
use AOI21X1  AOI21X1_401
timestamp 1696145522
transform -1 0 2796 0 -1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_68
timestamp 1696145522
transform -1 0 2820 0 -1 2105
box -2 -3 26 103
use AOI21X1  AOI21X1_33
timestamp 1696145522
transform -1 0 2852 0 -1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_69
timestamp 1696145522
transform 1 0 2852 0 -1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_915
timestamp 1696145522
transform -1 0 2908 0 -1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_399
timestamp 1696145522
transform -1 0 2940 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_914
timestamp 1696145522
transform -1 0 2972 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_919
timestamp 1696145522
transform -1 0 3004 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_918
timestamp 1696145522
transform -1 0 3036 0 -1 2105
box -2 -3 34 103
use FILL  FILL_20_5_0
timestamp 1696145522
transform 1 0 3036 0 -1 2105
box -2 -3 10 103
use FILL  FILL_20_5_1
timestamp 1696145522
transform 1 0 3044 0 -1 2105
box -2 -3 10 103
use AOI21X1  AOI21X1_395
timestamp 1696145522
transform 1 0 3052 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_910
timestamp 1696145522
transform 1 0 3084 0 -1 2105
box -2 -3 34 103
use NAND3X1  NAND3X1_54
timestamp 1696145522
transform -1 0 3148 0 -1 2105
box -2 -3 34 103
use XNOR2X1  XNOR2X1_28
timestamp 1696145522
transform -1 0 3204 0 -1 2105
box -2 -3 58 103
use NAND2X1  NAND2X1_83
timestamp 1696145522
transform -1 0 3228 0 -1 2105
box -2 -3 26 103
use NOR2X1  NOR2X1_120
timestamp 1696145522
transform 1 0 3228 0 -1 2105
box -2 -3 26 103
use INVX1  INVX1_33
timestamp 1696145522
transform -1 0 3268 0 -1 2105
box -2 -3 18 103
use XNOR2X1  XNOR2X1_29
timestamp 1696145522
transform -1 0 3324 0 -1 2105
box -2 -3 58 103
use BUFX4  BUFX4_104
timestamp 1696145522
transform 1 0 3324 0 -1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_920
timestamp 1696145522
transform -1 0 3388 0 -1 2105
box -2 -3 34 103
use INVX1  INVX1_322
timestamp 1696145522
transform -1 0 3404 0 -1 2105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_26
timestamp 1696145522
transform 1 0 3404 0 -1 2105
box -2 -3 98 103
use NOR2X1  NOR2X1_406
timestamp 1696145522
transform -1 0 3524 0 -1 2105
box -2 -3 26 103
use BUFX2  BUFX2_28
timestamp 1696145522
transform 1 0 3524 0 -1 2105
box -2 -3 26 103
use FILL  FILL_21_1
timestamp 1696145522
transform -1 0 3556 0 -1 2105
box -2 -3 10 103
use FILL  FILL_21_2
timestamp 1696145522
transform -1 0 3564 0 -1 2105
box -2 -3 10 103
use INVX1  INVX1_238
timestamp 1696145522
transform 1 0 4 0 1 2105
box -2 -3 18 103
use MUX2X1  MUX2X1_13
timestamp 1696145522
transform -1 0 68 0 1 2105
box -2 -3 50 103
use NAND2X1  NAND2X1_500
timestamp 1696145522
transform -1 0 92 0 1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_517
timestamp 1696145522
transform 1 0 92 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_577
timestamp 1696145522
transform -1 0 148 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_481
timestamp 1696145522
transform -1 0 172 0 1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_167
timestamp 1696145522
transform 1 0 172 0 1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_97
timestamp 1696145522
transform 1 0 196 0 1 2105
box -2 -3 26 103
use BUFX4  BUFX4_75
timestamp 1696145522
transform -1 0 252 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_454
timestamp 1696145522
transform 1 0 252 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_337
timestamp 1696145522
transform -1 0 308 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_294
timestamp 1696145522
transform 1 0 308 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_232
timestamp 1696145522
transform -1 0 364 0 1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_471
timestamp 1696145522
transform -1 0 388 0 1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_312
timestamp 1696145522
transform -1 0 412 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_457
timestamp 1696145522
transform -1 0 444 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_433
timestamp 1696145522
transform 1 0 444 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_405
timestamp 1696145522
transform -1 0 500 0 1 2105
box -2 -3 26 103
use FILL  FILL_21_0_0
timestamp 1696145522
transform 1 0 500 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_0_1
timestamp 1696145522
transform 1 0 508 0 1 2105
box -2 -3 10 103
use NAND2X1  NAND2X1_429
timestamp 1696145522
transform 1 0 516 0 1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_445
timestamp 1696145522
transform -1 0 564 0 1 2105
box -2 -3 26 103
use BUFX4  BUFX4_73
timestamp 1696145522
transform -1 0 596 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_391
timestamp 1696145522
transform -1 0 620 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_383
timestamp 1696145522
transform 1 0 620 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_357
timestamp 1696145522
transform 1 0 652 0 1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_378
timestamp 1696145522
transform -1 0 700 0 1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_208
timestamp 1696145522
transform 1 0 700 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_69
timestamp 1696145522
transform 1 0 724 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_120
timestamp 1696145522
transform 1 0 756 0 1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_209
timestamp 1696145522
transform -1 0 804 0 1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_123
timestamp 1696145522
transform 1 0 804 0 1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_152
timestamp 1696145522
transform 1 0 828 0 1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_249
timestamp 1696145522
transform -1 0 876 0 1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_259
timestamp 1696145522
transform 1 0 876 0 1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_174
timestamp 1696145522
transform -1 0 924 0 1 2105
box -2 -3 26 103
use BUFX4  BUFX4_71
timestamp 1696145522
transform -1 0 956 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_253
timestamp 1696145522
transform -1 0 980 0 1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_252
timestamp 1696145522
transform -1 0 1004 0 1 2105
box -2 -3 26 103
use FILL  FILL_21_1_0
timestamp 1696145522
transform -1 0 1012 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_1_1
timestamp 1696145522
transform -1 0 1020 0 1 2105
box -2 -3 10 103
use OAI21X1  OAI21X1_223
timestamp 1696145522
transform -1 0 1052 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_181
timestamp 1696145522
transform -1 0 1076 0 1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_179
timestamp 1696145522
transform -1 0 1100 0 1 2105
box -2 -3 26 103
use INVX1  INVX1_105
timestamp 1696145522
transform -1 0 1116 0 1 2105
box -2 -3 18 103
use NAND2X1  NAND2X1_413
timestamp 1696145522
transform 1 0 1116 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_440
timestamp 1696145522
transform -1 0 1172 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_127
timestamp 1696145522
transform 1 0 1172 0 1 2105
box -2 -3 26 103
use BUFX4  BUFX4_72
timestamp 1696145522
transform 1 0 1196 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_181
timestamp 1696145522
transform 1 0 1228 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_130
timestamp 1696145522
transform -1 0 1284 0 1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_214
timestamp 1696145522
transform -1 0 1308 0 1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_256
timestamp 1696145522
transform -1 0 1332 0 1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_588
timestamp 1696145522
transform 1 0 1332 0 1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_187
timestamp 1696145522
transform 1 0 1356 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_703
timestamp 1696145522
transform 1 0 1380 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_568
timestamp 1696145522
transform -1 0 1436 0 1 2105
box -2 -3 26 103
use MUX2X1  MUX2X1_78
timestamp 1696145522
transform 1 0 1436 0 1 2105
box -2 -3 50 103
use NOR2X1  NOR2X1_288
timestamp 1696145522
transform -1 0 1508 0 1 2105
box -2 -3 26 103
use FILL  FILL_21_2_0
timestamp 1696145522
transform -1 0 1516 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_2_1
timestamp 1696145522
transform -1 0 1524 0 1 2105
box -2 -3 10 103
use NAND3X1  NAND3X1_32
timestamp 1696145522
transform -1 0 1556 0 1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_362
timestamp 1696145522
transform -1 0 1580 0 1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_95
timestamp 1696145522
transform 1 0 1580 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_676
timestamp 1696145522
transform -1 0 1636 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_46
timestamp 1696145522
transform -1 0 1668 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_394
timestamp 1696145522
transform -1 0 1692 0 1 2105
box -2 -3 26 103
use INVX8  INVX8_13
timestamp 1696145522
transform 1 0 1692 0 1 2105
box -2 -3 42 103
use NAND2X1  NAND2X1_148
timestamp 1696145522
transform 1 0 1732 0 1 2105
box -2 -3 26 103
use BUFX4  BUFX4_5
timestamp 1696145522
transform -1 0 1788 0 1 2105
box -2 -3 34 103
use AND2X2  AND2X2_30
timestamp 1696145522
transform 1 0 1788 0 1 2105
box -2 -3 34 103
use AND2X2  AND2X2_31
timestamp 1696145522
transform 1 0 1820 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_445
timestamp 1696145522
transform 1 0 1852 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_451
timestamp 1696145522
transform 1 0 1884 0 1 2105
box -2 -3 34 103
use INVX1  INVX1_179
timestamp 1696145522
transform 1 0 1916 0 1 2105
box -2 -3 18 103
use NAND2X1  NAND2X1_408
timestamp 1696145522
transform -1 0 1956 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_450
timestamp 1696145522
transform 1 0 1956 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_407
timestamp 1696145522
transform 1 0 1988 0 1 2105
box -2 -3 26 103
use NOR2X1  NOR2X1_233
timestamp 1696145522
transform 1 0 2012 0 1 2105
box -2 -3 26 103
use FILL  FILL_21_3_0
timestamp 1696145522
transform -1 0 2044 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_3_1
timestamp 1696145522
transform -1 0 2052 0 1 2105
box -2 -3 10 103
use AOI21X1  AOI21X1_153
timestamp 1696145522
transform -1 0 2084 0 1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_232
timestamp 1696145522
transform -1 0 2108 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_474
timestamp 1696145522
transform -1 0 2140 0 1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_216
timestamp 1696145522
transform -1 0 2164 0 1 2105
box -2 -3 26 103
use AND2X2  AND2X2_21
timestamp 1696145522
transform 1 0 2164 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_438
timestamp 1696145522
transform 1 0 2196 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_461
timestamp 1696145522
transform 1 0 2228 0 1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_217
timestamp 1696145522
transform 1 0 2260 0 1 2105
box -2 -3 26 103
use AOI22X1  AOI22X1_13
timestamp 1696145522
transform -1 0 2324 0 1 2105
box -2 -3 42 103
use INVX4  INVX4_21
timestamp 1696145522
transform 1 0 2324 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_430
timestamp 1696145522
transform -1 0 2380 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_425
timestamp 1696145522
transform 1 0 2380 0 1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_226
timestamp 1696145522
transform 1 0 2412 0 1 2105
box -2 -3 26 103
use NOR2X1  NOR2X1_221
timestamp 1696145522
transform -1 0 2460 0 1 2105
box -2 -3 26 103
use AOI21X1  AOI21X1_145
timestamp 1696145522
transform 1 0 2460 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_238
timestamp 1696145522
transform 1 0 2492 0 1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_225
timestamp 1696145522
transform 1 0 2524 0 1 2105
box -2 -3 26 103
use FILL  FILL_21_4_0
timestamp 1696145522
transform -1 0 2556 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_4_1
timestamp 1696145522
transform -1 0 2564 0 1 2105
box -2 -3 10 103
use BUFX4  BUFX4_142
timestamp 1696145522
transform -1 0 2596 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_151
timestamp 1696145522
transform -1 0 2628 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_156
timestamp 1696145522
transform 1 0 2628 0 1 2105
box -2 -3 34 103
use AOI22X1  AOI22X1_55
timestamp 1696145522
transform 1 0 2660 0 1 2105
box -2 -3 42 103
use NOR2X1  NOR2X1_41
timestamp 1696145522
transform -1 0 2724 0 1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_52
timestamp 1696145522
transform -1 0 2748 0 1 2105
box -2 -3 26 103
use INVX4  INVX4_2
timestamp 1696145522
transform -1 0 2772 0 1 2105
box -2 -3 26 103
use AOI21X1  AOI21X1_16
timestamp 1696145522
transform 1 0 2772 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_912
timestamp 1696145522
transform -1 0 2836 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_913
timestamp 1696145522
transform -1 0 2868 0 1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_42
timestamp 1696145522
transform 1 0 2868 0 1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_57
timestamp 1696145522
transform 1 0 2892 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_652
timestamp 1696145522
transform -1 0 2948 0 1 2105
box -2 -3 34 103
use INVX1  INVX1_24
timestamp 1696145522
transform -1 0 2964 0 1 2105
box -2 -3 18 103
use NAND2X1  NAND2X1_59
timestamp 1696145522
transform 1 0 2964 0 1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_58
timestamp 1696145522
transform -1 0 3012 0 1 2105
box -2 -3 26 103
use NAND2X1  NAND2X1_56
timestamp 1696145522
transform -1 0 3036 0 1 2105
box -2 -3 26 103
use FILL  FILL_21_5_0
timestamp 1696145522
transform -1 0 3044 0 1 2105
box -2 -3 10 103
use FILL  FILL_21_5_1
timestamp 1696145522
transform -1 0 3052 0 1 2105
box -2 -3 10 103
use OAI21X1  OAI21X1_916
timestamp 1696145522
transform -1 0 3084 0 1 2105
box -2 -3 34 103
use XNOR2X1  XNOR2X1_47
timestamp 1696145522
transform 1 0 3084 0 1 2105
box -2 -3 58 103
use NAND3X1  NAND3X1_53
timestamp 1696145522
transform -1 0 3172 0 1 2105
box -2 -3 34 103
use BUFX4  BUFX4_141
timestamp 1696145522
transform -1 0 3204 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_167
timestamp 1696145522
transform -1 0 3236 0 1 2105
box -2 -3 34 103
use NAND2X1  NAND2X1_207
timestamp 1696145522
transform -1 0 3260 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_34
timestamp 1696145522
transform 1 0 3260 0 1 2105
box -2 -3 34 103
use AOI21X1  AOI21X1_60
timestamp 1696145522
transform -1 0 3324 0 1 2105
box -2 -3 34 103
use OAI21X1  OAI21X1_171
timestamp 1696145522
transform -1 0 3356 0 1 2105
box -2 -3 34 103
use NOR2X1  NOR2X1_70
timestamp 1696145522
transform -1 0 3380 0 1 2105
box -2 -3 26 103
use OAI21X1  OAI21X1_923
timestamp 1696145522
transform 1 0 3380 0 1 2105
box -2 -3 34 103
use AOI22X1  AOI22X1_1
timestamp 1696145522
transform 1 0 3412 0 1 2105
box -2 -3 42 103
use INVX1  INVX1_32
timestamp 1696145522
transform -1 0 3468 0 1 2105
box -2 -3 18 103
use INVX2  INVX2_31
timestamp 1696145522
transform -1 0 3484 0 1 2105
box -2 -3 18 103
use CLKBUF1  CLKBUF1_1
timestamp 1696145522
transform 1 0 3484 0 1 2105
box -2 -3 74 103
use FILL  FILL_22_1
timestamp 1696145522
transform 1 0 3556 0 1 2105
box -2 -3 10 103
use OAI21X1  OAI21X1_576
timestamp 1696145522
transform -1 0 36 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_112
timestamp 1696145522
transform 1 0 36 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_61
timestamp 1696145522
transform -1 0 92 0 -1 2305
box -2 -3 34 103
use MUX2X1  MUX2X1_59
timestamp 1696145522
transform -1 0 140 0 -1 2305
box -2 -3 50 103
use MUX2X1  MUX2X1_56
timestamp 1696145522
transform -1 0 188 0 -1 2305
box -2 -3 50 103
use MUX2X1  MUX2X1_53
timestamp 1696145522
transform -1 0 236 0 -1 2305
box -2 -3 50 103
use MUX2X1  MUX2X1_65
timestamp 1696145522
transform 1 0 236 0 -1 2305
box -2 -3 50 103
use OAI21X1  OAI21X1_258
timestamp 1696145522
transform -1 0 316 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_281
timestamp 1696145522
transform 1 0 316 0 -1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_386
timestamp 1696145522
transform 1 0 340 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_480
timestamp 1696145522
transform -1 0 396 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_422
timestamp 1696145522
transform -1 0 420 0 -1 2305
box -2 -3 26 103
use INVX1  INVX1_220
timestamp 1696145522
transform -1 0 436 0 -1 2305
box -2 -3 18 103
use OAI21X1  OAI21X1_526
timestamp 1696145522
transform -1 0 468 0 -1 2305
box -2 -3 34 103
use FILL  FILL_22_0_0
timestamp 1696145522
transform -1 0 476 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_0_1
timestamp 1696145522
transform -1 0 484 0 -1 2305
box -2 -3 10 103
use MUX2X1  MUX2X1_50
timestamp 1696145522
transform -1 0 532 0 -1 2305
box -2 -3 50 103
use OAI21X1  OAI21X1_432
timestamp 1696145522
transform -1 0 564 0 -1 2305
box -2 -3 34 103
use INVX1  INVX1_188
timestamp 1696145522
transform -1 0 580 0 -1 2305
box -2 -3 18 103
use INVX1  INVX1_130
timestamp 1696145522
transform -1 0 596 0 -1 2305
box -2 -3 18 103
use INVX1  INVX1_205
timestamp 1696145522
transform -1 0 612 0 -1 2305
box -2 -3 18 103
use MUX2X1  MUX2X1_10
timestamp 1696145522
transform 1 0 612 0 -1 2305
box -2 -3 50 103
use INVX1  INVX1_140
timestamp 1696145522
transform -1 0 676 0 -1 2305
box -2 -3 18 103
use OAI21X1  OAI21X1_456
timestamp 1696145522
transform 1 0 676 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_131
timestamp 1696145522
transform 1 0 708 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_80
timestamp 1696145522
transform -1 0 764 0 -1 2305
box -2 -3 34 103
use INVX1  INVX1_48
timestamp 1696145522
transform 1 0 764 0 -1 2305
box -2 -3 18 103
use INVX2  INVX2_46
timestamp 1696145522
transform 1 0 780 0 -1 2305
box -2 -3 18 103
use INVX1  INVX1_164
timestamp 1696145522
transform -1 0 812 0 -1 2305
box -2 -3 18 103
use MUX2X1  MUX2X1_8
timestamp 1696145522
transform -1 0 860 0 -1 2305
box -2 -3 50 103
use NAND2X1  NAND2X1_178
timestamp 1696145522
transform 1 0 860 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_412
timestamp 1696145522
transform -1 0 916 0 -1 2305
box -2 -3 34 103
use MUX2X1  MUX2X1_15
timestamp 1696145522
transform 1 0 916 0 -1 2305
box -2 -3 50 103
use MUX2X1  MUX2X1_18
timestamp 1696145522
transform -1 0 1012 0 -1 2305
box -2 -3 50 103
use FILL  FILL_22_1_0
timestamp 1696145522
transform -1 0 1020 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_1_1
timestamp 1696145522
transform -1 0 1028 0 -1 2305
box -2 -3 10 103
use OAI21X1  OAI21X1_467
timestamp 1696145522
transform -1 0 1060 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_137
timestamp 1696145522
transform -1 0 1092 0 -1 2305
box -2 -3 34 103
use INVX4  INVX4_14
timestamp 1696145522
transform 1 0 1092 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_275
timestamp 1696145522
transform -1 0 1148 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_142
timestamp 1696145522
transform -1 0 1180 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_217
timestamp 1696145522
transform 1 0 1180 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_106
timestamp 1696145522
transform -1 0 1244 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_151
timestamp 1696145522
transform -1 0 1268 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_143
timestamp 1696145522
transform 1 0 1268 0 -1 2305
box -2 -3 34 103
use MUX2X1  MUX2X1_77
timestamp 1696145522
transform -1 0 1348 0 -1 2305
box -2 -3 50 103
use NAND2X1  NAND2X1_96
timestamp 1696145522
transform 1 0 1348 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_47
timestamp 1696145522
transform -1 0 1404 0 -1 2305
box -2 -3 34 103
use MUX2X1  MUX2X1_68
timestamp 1696145522
transform -1 0 1452 0 -1 2305
box -2 -3 50 103
use NOR2X1  NOR2X1_208
timestamp 1696145522
transform 1 0 1452 0 -1 2305
box -2 -3 26 103
use INVX1  INVX1_173
timestamp 1696145522
transform 1 0 1476 0 -1 2305
box -2 -3 18 103
use NOR2X1  NOR2X1_209
timestamp 1696145522
transform -1 0 1516 0 -1 2305
box -2 -3 26 103
use FILL  FILL_22_2_0
timestamp 1696145522
transform 1 0 1516 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_2_1
timestamp 1696145522
transform 1 0 1524 0 -1 2305
box -2 -3 10 103
use NOR2X1  NOR2X1_210
timestamp 1696145522
transform 1 0 1532 0 -1 2305
box -2 -3 26 103
use INVX2  INVX2_74
timestamp 1696145522
transform -1 0 1572 0 -1 2305
box -2 -3 18 103
use OAI22X1  OAI22X1_7
timestamp 1696145522
transform -1 0 1612 0 -1 2305
box -2 -3 42 103
use AOI21X1  AOI21X1_134
timestamp 1696145522
transform -1 0 1644 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_551
timestamp 1696145522
transform 1 0 1644 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_669
timestamp 1696145522
transform -1 0 1700 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_552
timestamp 1696145522
transform -1 0 1724 0 -1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_425
timestamp 1696145522
transform 1 0 1724 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_464
timestamp 1696145522
transform 1 0 1748 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_427
timestamp 1696145522
transform 1 0 1780 0 -1 2305
box -2 -3 26 103
use INVX1  INVX1_194
timestamp 1696145522
transform 1 0 1804 0 -1 2305
box -2 -3 18 103
use AOI21X1  AOI21X1_164
timestamp 1696145522
transform 1 0 1820 0 -1 2305
box -2 -3 34 103
use AOI22X1  AOI22X1_17
timestamp 1696145522
transform 1 0 1852 0 -1 2305
box -2 -3 42 103
use INVX1  INVX1_185
timestamp 1696145522
transform 1 0 1892 0 -1 2305
box -2 -3 18 103
use XNOR2X1  XNOR2X1_35
timestamp 1696145522
transform -1 0 1964 0 -1 2305
box -2 -3 58 103
use NOR2X1  NOR2X1_231
timestamp 1696145522
transform 1 0 1964 0 -1 2305
box -2 -3 26 103
use AOI22X1  AOI22X1_16
timestamp 1696145522
transform 1 0 1988 0 -1 2305
box -2 -3 42 103
use FILL  FILL_22_3_0
timestamp 1696145522
transform -1 0 2036 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_3_1
timestamp 1696145522
transform -1 0 2044 0 -1 2305
box -2 -3 10 103
use OAI21X1  OAI21X1_454
timestamp 1696145522
transform -1 0 2076 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_452
timestamp 1696145522
transform -1 0 2108 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_421
timestamp 1696145522
transform -1 0 2132 0 -1 2305
box -2 -3 26 103
use AOI21X1  AOI21X1_162
timestamp 1696145522
transform 1 0 2132 0 -1 2305
box -2 -3 34 103
use INVX2  INVX2_75
timestamp 1696145522
transform 1 0 2164 0 -1 2305
box -2 -3 18 103
use NOR2X1  NOR2X1_220
timestamp 1696145522
transform 1 0 2180 0 -1 2305
box -2 -3 26 103
use INVX1  INVX1_186
timestamp 1696145522
transform 1 0 2204 0 -1 2305
box -2 -3 18 103
use OR2X2  OR2X2_24
timestamp 1696145522
transform 1 0 2220 0 -1 2305
box -2 -3 34 103
use AND2X2  AND2X2_24
timestamp 1696145522
transform 1 0 2252 0 -1 2305
box -2 -3 34 103
use BUFX4  BUFX4_57
timestamp 1696145522
transform -1 0 2316 0 -1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_234
timestamp 1696145522
transform -1 0 2340 0 -1 2305
box -2 -3 26 103
use AOI21X1  AOI21X1_157
timestamp 1696145522
transform 1 0 2340 0 -1 2305
box -2 -3 34 103
use INVX4  INVX4_16
timestamp 1696145522
transform -1 0 2396 0 -1 2305
box -2 -3 26 103
use AOI22X1  AOI22X1_5
timestamp 1696145522
transform 1 0 2396 0 -1 2305
box -2 -3 42 103
use NAND2X1  NAND2X1_237
timestamp 1696145522
transform -1 0 2460 0 -1 2305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_46
timestamp 1696145522
transform 1 0 2460 0 -1 2305
box -2 -3 98 103
use FILL  FILL_22_4_0
timestamp 1696145522
transform 1 0 2556 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_4_1
timestamp 1696145522
transform 1 0 2564 0 -1 2305
box -2 -3 10 103
use AOI21X1  AOI21X1_68
timestamp 1696145522
transform 1 0 2572 0 -1 2305
box -2 -3 34 103
use BUFX4  BUFX4_6
timestamp 1696145522
transform 1 0 2604 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_649
timestamp 1696145522
transform -1 0 2660 0 -1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_503
timestamp 1696145522
transform -1 0 2684 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_935
timestamp 1696145522
transform 1 0 2684 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_648
timestamp 1696145522
transform -1 0 2740 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_934
timestamp 1696145522
transform -1 0 2772 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_646
timestamp 1696145522
transform -1 0 2796 0 -1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_500
timestamp 1696145522
transform 1 0 2796 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_929
timestamp 1696145522
transform -1 0 2852 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_928
timestamp 1696145522
transform 1 0 2852 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_927
timestamp 1696145522
transform -1 0 2916 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_921
timestamp 1696145522
transform -1 0 2948 0 -1 2305
box -2 -3 34 103
use XNOR2X1  XNOR2X1_27
timestamp 1696145522
transform -1 0 3004 0 -1 2305
box -2 -3 58 103
use OAI21X1  OAI21X1_22
timestamp 1696145522
transform 1 0 3004 0 -1 2305
box -2 -3 34 103
use FILL  FILL_22_5_0
timestamp 1696145522
transform 1 0 3036 0 -1 2305
box -2 -3 10 103
use FILL  FILL_22_5_1
timestamp 1696145522
transform 1 0 3044 0 -1 2305
box -2 -3 10 103
use OAI21X1  OAI21X1_21
timestamp 1696145522
transform 1 0 3052 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_20
timestamp 1696145522
transform -1 0 3116 0 -1 2305
box -2 -3 34 103
use INVX2  INVX2_29
timestamp 1696145522
transform 1 0 3116 0 -1 2305
box -2 -3 18 103
use NAND2X1  NAND2X1_46
timestamp 1696145522
transform 1 0 3132 0 -1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_45
timestamp 1696145522
transform 1 0 3156 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_170
timestamp 1696145522
transform 1 0 3180 0 -1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_33
timestamp 1696145522
transform 1 0 3212 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_647
timestamp 1696145522
transform 1 0 3244 0 -1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_932
timestamp 1696145522
transform -1 0 3300 0 -1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_49
timestamp 1696145522
transform 1 0 3300 0 -1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_50
timestamp 1696145522
transform -1 0 3348 0 -1 2305
box -2 -3 26 103
use INVX1  INVX1_325
timestamp 1696145522
transform 1 0 3348 0 -1 2305
box -2 -3 18 103
use OAI21X1  OAI21X1_930
timestamp 1696145522
transform 1 0 3364 0 -1 2305
box -2 -3 34 103
use INVX1  INVX1_22
timestamp 1696145522
transform 1 0 3396 0 -1 2305
box -2 -3 18 103
use NAND2X1  NAND2X1_48
timestamp 1696145522
transform -1 0 3436 0 -1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_44
timestamp 1696145522
transform -1 0 3460 0 -1 2305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_28
timestamp 1696145522
transform 1 0 3460 0 -1 2305
box -2 -3 98 103
use FILL  FILL_23_1
timestamp 1696145522
transform -1 0 3564 0 -1 2305
box -2 -3 10 103
use NAND2X1  NAND2X1_499
timestamp 1696145522
transform -1 0 28 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_126
timestamp 1696145522
transform 1 0 28 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_604
timestamp 1696145522
transform -1 0 92 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_586
timestamp 1696145522
transform 1 0 92 0 1 2305
box -2 -3 34 103
use MUX2X1  MUX2X1_5
timestamp 1696145522
transform 1 0 124 0 1 2305
box -2 -3 50 103
use OAI21X1  OAI21X1_64
timestamp 1696145522
transform -1 0 204 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_567
timestamp 1696145522
transform 1 0 204 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_372
timestamp 1696145522
transform -1 0 268 0 1 2305
box -2 -3 34 103
use INVX1  INVX1_159
timestamp 1696145522
transform -1 0 284 0 1 2305
box -2 -3 18 103
use NAND2X1  NAND2X1_348
timestamp 1696145522
transform -1 0 308 0 1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_369
timestamp 1696145522
transform 1 0 308 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_401
timestamp 1696145522
transform 1 0 332 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_439
timestamp 1696145522
transform -1 0 388 0 1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_114
timestamp 1696145522
transform 1 0 388 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_504
timestamp 1696145522
transform 1 0 412 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_451
timestamp 1696145522
transform 1 0 444 0 1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_466
timestamp 1696145522
transform 1 0 468 0 1 2305
box -2 -3 26 103
use FILL  FILL_23_0_0
timestamp 1696145522
transform -1 0 500 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_0_1
timestamp 1696145522
transform -1 0 508 0 1 2305
box -2 -3 10 103
use INVX1  INVX1_171
timestamp 1696145522
transform -1 0 524 0 1 2305
box -2 -3 18 103
use NAND2X1  NAND2X1_404
timestamp 1696145522
transform 1 0 524 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_63
timestamp 1696145522
transform -1 0 580 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_547
timestamp 1696145522
transform 1 0 580 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_122
timestamp 1696145522
transform 1 0 612 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_479
timestamp 1696145522
transform -1 0 668 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_71
timestamp 1696145522
transform -1 0 700 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_491
timestamp 1696145522
transform -1 0 732 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_444
timestamp 1696145522
transform 1 0 732 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_70
timestamp 1696145522
transform -1 0 788 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_371
timestamp 1696145522
transform -1 0 820 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_129
timestamp 1696145522
transform 1 0 820 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_382
timestamp 1696145522
transform -1 0 884 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_135
timestamp 1696145522
transform -1 0 916 0 1 2305
box -2 -3 34 103
use INVX2  INVX2_73
timestamp 1696145522
transform -1 0 932 0 1 2305
box -2 -3 18 103
use AND2X2  AND2X2_40
timestamp 1696145522
transform 1 0 932 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_82
timestamp 1696145522
transform 1 0 964 0 1 2305
box -2 -3 34 103
use FILL  FILL_23_1_0
timestamp 1696145522
transform 1 0 996 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_1_1
timestamp 1696145522
transform 1 0 1004 0 1 2305
box -2 -3 10 103
use NAND2X1  NAND2X1_180
timestamp 1696145522
transform 1 0 1012 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_322
timestamp 1696145522
transform 1 0 1036 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_335
timestamp 1696145522
transform -1 0 1092 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_140
timestamp 1696145522
transform -1 0 1124 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_185
timestamp 1696145522
transform 1 0 1124 0 1 2305
box -2 -3 26 103
use MUX2X1  MUX2X1_6
timestamp 1696145522
transform 1 0 1148 0 1 2305
box -2 -3 50 103
use NAND2X1  NAND2X1_311
timestamp 1696145522
transform 1 0 1196 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_293
timestamp 1696145522
transform -1 0 1252 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_75
timestamp 1696145522
transform 1 0 1252 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_186
timestamp 1696145522
transform 1 0 1284 0 1 2305
box -2 -3 26 103
use INVX2  INVX2_43
timestamp 1696145522
transform 1 0 1308 0 1 2305
box -2 -3 18 103
use NAND3X1  NAND3X1_41
timestamp 1696145522
transform -1 0 1356 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_150
timestamp 1696145522
transform 1 0 1356 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_105
timestamp 1696145522
transform -1 0 1412 0 1 2305
box -2 -3 34 103
use BUFX4  BUFX4_4
timestamp 1696145522
transform -1 0 1444 0 1 2305
box -2 -3 34 103
use INVX1  INVX1_190
timestamp 1696145522
transform -1 0 1460 0 1 2305
box -2 -3 18 103
use OAI21X1  OAI21X1_671
timestamp 1696145522
transform 1 0 1460 0 1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_292
timestamp 1696145522
transform 1 0 1492 0 1 2305
box -2 -3 34 103
use FILL  FILL_23_2_0
timestamp 1696145522
transform 1 0 1524 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_2_1
timestamp 1696145522
transform 1 0 1532 0 1 2305
box -2 -3 10 103
use AOI21X1  AOI21X1_140
timestamp 1696145522
transform 1 0 1540 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_426
timestamp 1696145522
transform 1 0 1572 0 1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_438
timestamp 1696145522
transform 1 0 1596 0 1 2305
box -2 -3 26 103
use INVX1  INVX1_191
timestamp 1696145522
transform -1 0 1636 0 1 2305
box -2 -3 18 103
use NOR2X1  NOR2X1_250
timestamp 1696145522
transform -1 0 1660 0 1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_423
timestamp 1696145522
transform -1 0 1684 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_673
timestamp 1696145522
transform 1 0 1684 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_668
timestamp 1696145522
transform -1 0 1748 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_476
timestamp 1696145522
transform -1 0 1780 0 1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_422
timestamp 1696145522
transform 1 0 1780 0 1 2305
box -2 -3 26 103
use OR2X2  OR2X2_29
timestamp 1696145522
transform -1 0 1836 0 1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_264
timestamp 1696145522
transform 1 0 1836 0 1 2305
box -2 -3 26 103
use OR2X2  OR2X2_30
timestamp 1696145522
transform 1 0 1860 0 1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_249
timestamp 1696145522
transform 1 0 1892 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_475
timestamp 1696145522
transform -1 0 1948 0 1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_230
timestamp 1696145522
transform 1 0 1948 0 1 2305
box -2 -3 26 103
use INVX1  INVX1_184
timestamp 1696145522
transform -1 0 1988 0 1 2305
box -2 -3 18 103
use NOR2X1  NOR2X1_229
timestamp 1696145522
transform -1 0 2012 0 1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_238
timestamp 1696145522
transform -1 0 2036 0 1 2305
box -2 -3 26 103
use FILL  FILL_23_3_0
timestamp 1696145522
transform -1 0 2044 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_3_1
timestamp 1696145522
transform -1 0 2052 0 1 2305
box -2 -3 10 103
use NAND3X1  NAND3X1_29
timestamp 1696145522
transform -1 0 2084 0 1 2305
box -2 -3 34 103
use OR2X2  OR2X2_28
timestamp 1696145522
transform -1 0 2116 0 1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_244
timestamp 1696145522
transform 1 0 2116 0 1 2305
box -2 -3 26 103
use NAND2X1  NAND2X1_432
timestamp 1696145522
transform -1 0 2164 0 1 2305
box -2 -3 26 103
use AOI21X1  AOI21X1_159
timestamp 1696145522
transform -1 0 2196 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_410
timestamp 1696145522
transform -1 0 2220 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_462
timestamp 1696145522
transform 1 0 2220 0 1 2305
box -2 -3 34 103
use INVX4  INVX4_22
timestamp 1696145522
transform -1 0 2276 0 1 2305
box -2 -3 26 103
use NAND3X1  NAND3X1_26
timestamp 1696145522
transform 1 0 2276 0 1 2305
box -2 -3 34 103
use INVX1  INVX1_192
timestamp 1696145522
transform -1 0 2324 0 1 2305
box -2 -3 18 103
use OAI21X1  OAI21X1_463
timestamp 1696145522
transform 1 0 2324 0 1 2305
box -2 -3 34 103
use NAND3X1  NAND3X1_27
timestamp 1696145522
transform -1 0 2388 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_598
timestamp 1696145522
transform -1 0 2420 0 1 2305
box -2 -3 34 103
use XNOR2X1  XNOR2X1_30
timestamp 1696145522
transform -1 0 2476 0 1 2305
box -2 -3 58 103
use OAI21X1  OAI21X1_205
timestamp 1696145522
transform 1 0 2476 0 1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_64
timestamp 1696145522
transform -1 0 2540 0 1 2305
box -2 -3 34 103
use FILL  FILL_23_4_0
timestamp 1696145522
transform -1 0 2548 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_4_1
timestamp 1696145522
transform -1 0 2556 0 1 2305
box -2 -3 10 103
use AOI21X1  AOI21X1_62
timestamp 1696145522
transform -1 0 2588 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_169
timestamp 1696145522
transform -1 0 2620 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_202
timestamp 1696145522
transform 1 0 2620 0 1 2305
box -2 -3 34 103
use AOI22X1  AOI22X1_4
timestamp 1696145522
transform -1 0 2692 0 1 2305
box -2 -3 42 103
use BUFX4  BUFX4_63
timestamp 1696145522
transform 1 0 2692 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_154
timestamp 1696145522
transform 1 0 2724 0 1 2305
box -2 -3 34 103
use XNOR2X1  XNOR2X1_26
timestamp 1696145522
transform 1 0 2756 0 1 2305
box -2 -3 58 103
use OAI21X1  OAI21X1_936
timestamp 1696145522
transform -1 0 2844 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_82
timestamp 1696145522
transform 1 0 2844 0 1 2305
box -2 -3 26 103
use AOI21X1  AOI21X1_47
timestamp 1696145522
transform -1 0 2900 0 1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_106
timestamp 1696145522
transform -1 0 2924 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_151
timestamp 1696145522
transform 1 0 2924 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_192
timestamp 1696145522
transform -1 0 2980 0 1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_104
timestamp 1696145522
transform -1 0 3004 0 1 2305
box -2 -3 26 103
use OR2X2  OR2X2_2
timestamp 1696145522
transform 1 0 3004 0 1 2305
box -2 -3 34 103
use NOR2X1  NOR2X1_110
timestamp 1696145522
transform -1 0 3060 0 1 2305
box -2 -3 26 103
use FILL  FILL_23_5_0
timestamp 1696145522
transform -1 0 3068 0 1 2305
box -2 -3 10 103
use FILL  FILL_23_5_1
timestamp 1696145522
transform -1 0 3076 0 1 2305
box -2 -3 10 103
use OAI21X1  OAI21X1_23
timestamp 1696145522
transform -1 0 3108 0 1 2305
box -2 -3 34 103
use INVX2  INVX2_2
timestamp 1696145522
transform 1 0 3108 0 1 2305
box -2 -3 18 103
use AOI21X1  AOI21X1_286
timestamp 1696145522
transform -1 0 3156 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_47
timestamp 1696145522
transform -1 0 3180 0 1 2305
box -2 -3 26 103
use OAI21X1  OAI21X1_653
timestamp 1696145522
transform -1 0 3212 0 1 2305
box -2 -3 34 103
use NAND2X1  NAND2X1_51
timestamp 1696145522
transform 1 0 3212 0 1 2305
box -2 -3 26 103
use NOR2X1  NOR2X1_67
timestamp 1696145522
transform 1 0 3236 0 1 2305
box -2 -3 26 103
use XNOR2X1  XNOR2X1_48
timestamp 1696145522
transform 1 0 3260 0 1 2305
box -2 -3 58 103
use AOI21X1  AOI21X1_407
timestamp 1696145522
transform -1 0 3348 0 1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_402
timestamp 1696145522
transform 1 0 3348 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_922
timestamp 1696145522
transform 1 0 3380 0 1 2305
box -2 -3 34 103
use AOI21X1  AOI21X1_405
timestamp 1696145522
transform 1 0 3412 0 1 2305
box -2 -3 34 103
use OAI21X1  OAI21X1_931
timestamp 1696145522
transform 1 0 3444 0 1 2305
box -2 -3 34 103
use AOI22X1  AOI22X1_57
timestamp 1696145522
transform -1 0 3516 0 1 2305
box -2 -3 42 103
use INVX1  INVX1_274
timestamp 1696145522
transform -1 0 3532 0 1 2305
box -2 -3 18 103
use BUFX2  BUFX2_30
timestamp 1696145522
transform 1 0 3532 0 1 2305
box -2 -3 26 103
use FILL  FILL_24_1
timestamp 1696145522
transform 1 0 3556 0 1 2305
box -2 -3 10 103
use OAI21X1  OAI21X1_591
timestamp 1696145522
transform 1 0 4 0 -1 2505
box -2 -3 34 103
use INVX4  INVX4_12
timestamp 1696145522
transform -1 0 60 0 -1 2505
box -2 -3 26 103
use INVX2  INVX2_87
timestamp 1696145522
transform 1 0 60 0 -1 2505
box -2 -3 18 103
use NAND2X1  NAND2X1_115
timestamp 1696145522
transform 1 0 76 0 -1 2505
box -2 -3 26 103
use OAI22X1  OAI22X1_24
timestamp 1696145522
transform 1 0 100 0 -1 2505
box -2 -3 42 103
use INVX1  INVX1_252
timestamp 1696145522
transform 1 0 140 0 -1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_656
timestamp 1696145522
transform -1 0 188 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_354
timestamp 1696145522
transform -1 0 212 0 -1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_355
timestamp 1696145522
transform -1 0 236 0 -1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_522
timestamp 1696145522
transform -1 0 260 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_624
timestamp 1696145522
transform -1 0 292 0 -1 2505
box -2 -3 34 103
use AOI22X1  AOI22X1_28
timestamp 1696145522
transform 1 0 292 0 -1 2505
box -2 -3 42 103
use INVX1  INVX1_255
timestamp 1696145522
transform -1 0 348 0 -1 2505
box -2 -3 18 103
use INVX4  INVX4_10
timestamp 1696145522
transform -1 0 372 0 -1 2505
box -2 -3 26 103
use MUX2X1  MUX2X1_14
timestamp 1696145522
transform -1 0 420 0 -1 2505
box -2 -3 50 103
use OAI21X1  OAI21X1_617
timestamp 1696145522
transform -1 0 452 0 -1 2505
box -2 -3 34 103
use INVX1  INVX1_97
timestamp 1696145522
transform -1 0 468 0 -1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_534
timestamp 1696145522
transform -1 0 500 0 -1 2505
box -2 -3 34 103
use FILL  FILL_24_0_0
timestamp 1696145522
transform 1 0 500 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_0_1
timestamp 1696145522
transform 1 0 508 0 -1 2505
box -2 -3 10 103
use NAND2X1  NAND2X1_470
timestamp 1696145522
transform 1 0 516 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_556
timestamp 1696145522
transform -1 0 572 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_131
timestamp 1696145522
transform -1 0 604 0 -1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_118
timestamp 1696145522
transform -1 0 628 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_67
timestamp 1696145522
transform -1 0 660 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_525
timestamp 1696145522
transform 1 0 660 0 -1 2505
box -2 -3 34 103
use INVX1  INVX1_210
timestamp 1696145522
transform -1 0 708 0 -1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_503
timestamp 1696145522
transform -1 0 740 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_68
timestamp 1696145522
transform 1 0 740 0 -1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_119
timestamp 1696145522
transform 1 0 772 0 -1 2505
box -2 -3 26 103
use MUX2X1  MUX2X1_16
timestamp 1696145522
transform -1 0 844 0 -1 2505
box -2 -3 50 103
use OAI21X1  OAI21X1_511
timestamp 1696145522
transform -1 0 876 0 -1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_377
timestamp 1696145522
transform 1 0 876 0 -1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_368
timestamp 1696145522
transform 1 0 900 0 -1 2505
box -2 -3 26 103
use MUX2X1  MUX2X1_17
timestamp 1696145522
transform 1 0 924 0 -1 2505
box -2 -3 50 103
use OAI21X1  OAI21X1_400
timestamp 1696145522
transform -1 0 1004 0 -1 2505
box -2 -3 34 103
use FILL  FILL_24_1_0
timestamp 1696145522
transform -1 0 1012 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_1_1
timestamp 1696145522
transform -1 0 1020 0 -1 2505
box -2 -3 10 103
use MUX2X1  MUX2X1_9
timestamp 1696145522
transform -1 0 1068 0 -1 2505
box -2 -3 50 103
use NAND2X1  NAND2X1_183
timestamp 1696145522
transform 1 0 1068 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_348
timestamp 1696145522
transform -1 0 1124 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_257
timestamp 1696145522
transform -1 0 1156 0 -1 2505
box -2 -3 34 103
use MUX2X1  MUX2X1_19
timestamp 1696145522
transform -1 0 1204 0 -1 2505
box -2 -3 50 103
use NAND2X1  NAND2X1_129
timestamp 1696145522
transform 1 0 1204 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_77
timestamp 1696145522
transform -1 0 1260 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_336
timestamp 1696145522
transform -1 0 1292 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_198
timestamp 1696145522
transform 1 0 1292 0 -1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_231
timestamp 1696145522
transform -1 0 1348 0 -1 2505
box -2 -3 26 103
use MUX2X1  MUX2X1_7
timestamp 1696145522
transform -1 0 1396 0 -1 2505
box -2 -3 50 103
use INVX2  INVX2_45
timestamp 1696145522
transform 1 0 1396 0 -1 2505
box -2 -3 18 103
use INVX2  INVX2_56
timestamp 1696145522
transform 1 0 1412 0 -1 2505
box -2 -3 18 103
use BUFX4  BUFX4_58
timestamp 1696145522
transform 1 0 1428 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_670
timestamp 1696145522
transform 1 0 1460 0 -1 2505
box -2 -3 34 103
use NAND3X1  NAND3X1_21
timestamp 1696145522
transform 1 0 1492 0 -1 2505
box -2 -3 34 103
use FILL  FILL_24_2_0
timestamp 1696145522
transform -1 0 1532 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_2_1
timestamp 1696145522
transform -1 0 1540 0 -1 2505
box -2 -3 10 103
use NAND2X1  NAND2X1_398
timestamp 1696145522
transform -1 0 1564 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_421
timestamp 1696145522
transform 1 0 1564 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_200
timestamp 1696145522
transform -1 0 1620 0 -1 2505
box -2 -3 26 103
use BUFX4  BUFX4_157
timestamp 1696145522
transform -1 0 1652 0 -1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_133
timestamp 1696145522
transform 1 0 1652 0 -1 2505
box -2 -3 34 103
use OR2X2  OR2X2_21
timestamp 1696145522
transform 1 0 1684 0 -1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_136
timestamp 1696145522
transform 1 0 1716 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_424
timestamp 1696145522
transform -1 0 1780 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_247
timestamp 1696145522
transform -1 0 1804 0 -1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_219
timestamp 1696145522
transform -1 0 1828 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_499
timestamp 1696145522
transform 1 0 1828 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_248
timestamp 1696145522
transform 1 0 1860 0 -1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_251
timestamp 1696145522
transform -1 0 1908 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_422
timestamp 1696145522
transform -1 0 1940 0 -1 2505
box -2 -3 34 103
use INVX1  INVX1_200
timestamp 1696145522
transform 1 0 1940 0 -1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_477
timestamp 1696145522
transform -1 0 1988 0 -1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_166
timestamp 1696145522
transform -1 0 2020 0 -1 2505
box -2 -3 34 103
use FILL  FILL_24_3_0
timestamp 1696145522
transform -1 0 2028 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_3_1
timestamp 1696145522
transform -1 0 2036 0 -1 2505
box -2 -3 10 103
use INVX1  INVX1_199
timestamp 1696145522
transform -1 0 2052 0 -1 2505
box -2 -3 18 103
use AOI21X1  AOI21X1_113
timestamp 1696145522
transform 1 0 2052 0 -1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_434
timestamp 1696145522
transform 1 0 2084 0 -1 2505
box -2 -3 26 103
use AOI21X1  AOI21X1_141
timestamp 1696145522
transform -1 0 2140 0 -1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_433
timestamp 1696145522
transform 1 0 2140 0 -1 2505
box -2 -3 26 103
use BUFX4  BUFX4_139
timestamp 1696145522
transform -1 0 2196 0 -1 2505
box -2 -3 34 103
use BUFX4  BUFX4_143
timestamp 1696145522
transform -1 0 2228 0 -1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_152
timestamp 1696145522
transform 1 0 2228 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_453
timestamp 1696145522
transform 1 0 2260 0 -1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_322
timestamp 1696145522
transform -1 0 2316 0 -1 2505
box -2 -3 26 103
use AOI21X1  AOI21X1_139
timestamp 1696145522
transform 1 0 2316 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_423
timestamp 1696145522
transform 1 0 2348 0 -1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_163
timestamp 1696145522
transform 1 0 2380 0 -1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_549
timestamp 1696145522
transform -1 0 2436 0 -1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_138
timestamp 1696145522
transform -1 0 2460 0 -1 2505
box -2 -3 26 103
use AOI21X1  AOI21X1_70
timestamp 1696145522
transform -1 0 2492 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_137
timestamp 1696145522
transform -1 0 2516 0 -1 2505
box -2 -3 26 103
use OR2X2  OR2X2_6
timestamp 1696145522
transform 1 0 2516 0 -1 2505
box -2 -3 34 103
use FILL  FILL_24_4_0
timestamp 1696145522
transform 1 0 2548 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_4_1
timestamp 1696145522
transform 1 0 2556 0 -1 2505
box -2 -3 10 103
use AOI21X1  AOI21X1_146
timestamp 1696145522
transform 1 0 2564 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_242
timestamp 1696145522
transform -1 0 2628 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_102
timestamp 1696145522
transform 1 0 2628 0 -1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_103
timestamp 1696145522
transform 1 0 2652 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_239
timestamp 1696145522
transform -1 0 2708 0 -1 2505
box -2 -3 34 103
use INVX4  INVX4_15
timestamp 1696145522
transform 1 0 2708 0 -1 2505
box -2 -3 26 103
use NAND3X1  NAND3X1_5
timestamp 1696145522
transform 1 0 2732 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_204
timestamp 1696145522
transform 1 0 2764 0 -1 2505
box -2 -3 34 103
use NAND3X1  NAND3X1_6
timestamp 1696145522
transform -1 0 2828 0 -1 2505
box -2 -3 34 103
use BUFX4  BUFX4_158
timestamp 1696145522
transform 1 0 2828 0 -1 2505
box -2 -3 34 103
use INVX8  INVX8_6
timestamp 1696145522
transform 1 0 2860 0 -1 2505
box -2 -3 42 103
use BUFX4  BUFX4_99
timestamp 1696145522
transform 1 0 2900 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_942
timestamp 1696145522
transform 1 0 2932 0 -1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_650
timestamp 1696145522
transform -1 0 2988 0 -1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_505
timestamp 1696145522
transform 1 0 2988 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_941
timestamp 1696145522
transform 1 0 3012 0 -1 2505
box -2 -3 34 103
use FILL  FILL_24_5_0
timestamp 1696145522
transform 1 0 3044 0 -1 2505
box -2 -3 10 103
use FILL  FILL_24_5_1
timestamp 1696145522
transform 1 0 3052 0 -1 2505
box -2 -3 10 103
use INVX1  INVX1_25
timestamp 1696145522
transform 1 0 3060 0 -1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_940
timestamp 1696145522
transform -1 0 3108 0 -1 2505
box -2 -3 34 103
use INVX1  INVX1_327
timestamp 1696145522
transform -1 0 3124 0 -1 2505
box -2 -3 18 103
use NAND2X1  NAND2X1_540
timestamp 1696145522
transform 1 0 3124 0 -1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_506
timestamp 1696145522
transform -1 0 3172 0 -1 2505
box -2 -3 26 103
use AOI21X1  AOI21X1_408
timestamp 1696145522
transform 1 0 3172 0 -1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_938
timestamp 1696145522
transform -1 0 3236 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_121
timestamp 1696145522
transform 1 0 3236 0 -1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_651
timestamp 1696145522
transform 1 0 3260 0 -1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_944
timestamp 1696145522
transform -1 0 3316 0 -1 2505
box -2 -3 34 103
use XNOR2X1  XNOR2X1_49
timestamp 1696145522
transform 1 0 3316 0 -1 2505
box -2 -3 58 103
use OAI21X1  OAI21X1_924
timestamp 1696145522
transform -1 0 3404 0 -1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_403
timestamp 1696145522
transform 1 0 3404 0 -1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_501
timestamp 1696145522
transform 1 0 3436 0 -1 2505
box -2 -3 26 103
use AOI22X1  AOI22X1_56
timestamp 1696145522
transform -1 0 3500 0 -1 2505
box -2 -3 42 103
use INVX1  INVX1_275
timestamp 1696145522
transform -1 0 3516 0 -1 2505
box -2 -3 18 103
use NAND3X1  NAND3X1_50
timestamp 1696145522
transform 1 0 3516 0 -1 2505
box -2 -3 34 103
use FILL  FILL_25_1
timestamp 1696145522
transform -1 0 3556 0 -1 2505
box -2 -3 10 103
use FILL  FILL_25_2
timestamp 1696145522
transform -1 0 3564 0 -1 2505
box -2 -3 10 103
use INVX4  INVX4_9
timestamp 1696145522
transform 1 0 4 0 1 2505
box -2 -3 26 103
use INVX4  INVX4_13
timestamp 1696145522
transform 1 0 28 0 1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_170
timestamp 1696145522
transform -1 0 76 0 1 2505
box -2 -3 26 103
use INVX1  INVX1_245
timestamp 1696145522
transform 1 0 76 0 1 2505
box -2 -3 18 103
use NOR2X1  NOR2X1_343
timestamp 1696145522
transform -1 0 116 0 1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_358
timestamp 1696145522
transform -1 0 140 0 1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_342
timestamp 1696145522
transform -1 0 164 0 1 2505
box -2 -3 26 103
use INVX2  INVX2_39
timestamp 1696145522
transform 1 0 164 0 1 2505
box -2 -3 18 103
use AND2X2  AND2X2_39
timestamp 1696145522
transform 1 0 180 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_622
timestamp 1696145522
transform 1 0 212 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_612
timestamp 1696145522
transform -1 0 276 0 1 2505
box -2 -3 34 103
use INVX2  INVX2_90
timestamp 1696145522
transform 1 0 276 0 1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_571
timestamp 1696145522
transform 1 0 292 0 1 2505
box -2 -3 34 103
use AND2X2  AND2X2_37
timestamp 1696145522
transform 1 0 324 0 1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_344
timestamp 1696145522
transform -1 0 380 0 1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_359
timestamp 1696145522
transform 1 0 380 0 1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_350
timestamp 1696145522
transform 1 0 404 0 1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_351
timestamp 1696145522
transform 1 0 428 0 1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_602
timestamp 1696145522
transform -1 0 484 0 1 2505
box -2 -3 34 103
use FILL  FILL_25_0_0
timestamp 1696145522
transform -1 0 492 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_0_1
timestamp 1696145522
transform -1 0 500 0 1 2505
box -2 -3 10 103
use AOI21X1  AOI21X1_252
timestamp 1696145522
transform -1 0 532 0 1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_289
timestamp 1696145522
transform 1 0 532 0 1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_175
timestamp 1696145522
transform 1 0 564 0 1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_352
timestamp 1696145522
transform -1 0 612 0 1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_364
timestamp 1696145522
transform -1 0 636 0 1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_526
timestamp 1696145522
transform 1 0 636 0 1 2505
box -2 -3 26 103
use INVX1  INVX1_256
timestamp 1696145522
transform -1 0 676 0 1 2505
box -2 -3 18 103
use NOR2X1  NOR2X1_365
timestamp 1696145522
transform -1 0 700 0 1 2505
box -2 -3 26 103
use NAND3X1  NAND3X1_55
timestamp 1696145522
transform 1 0 700 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_637
timestamp 1696145522
transform -1 0 764 0 1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_121
timestamp 1696145522
transform 1 0 764 0 1 2505
box -2 -3 26 103
use INVX4  INVX4_25
timestamp 1696145522
transform -1 0 812 0 1 2505
box -2 -3 26 103
use NAND3X1  NAND3X1_40
timestamp 1696145522
transform -1 0 844 0 1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_173
timestamp 1696145522
transform 1 0 844 0 1 2505
box -2 -3 26 103
use INVX1  INVX1_211
timestamp 1696145522
transform 1 0 868 0 1 2505
box -2 -3 18 103
use INVX2  INVX2_47
timestamp 1696145522
transform -1 0 900 0 1 2505
box -2 -3 18 103
use NAND2X1  NAND2X1_523
timestamp 1696145522
transform -1 0 924 0 1 2505
box -2 -3 26 103
use AND2X2  AND2X2_34
timestamp 1696145522
transform 1 0 924 0 1 2505
box -2 -3 34 103
use AND2X2  AND2X2_42
timestamp 1696145522
transform 1 0 956 0 1 2505
box -2 -3 34 103
use FILL  FILL_25_1_0
timestamp 1696145522
transform 1 0 988 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_1_1
timestamp 1696145522
transform 1 0 996 0 1 2505
box -2 -3 10 103
use AND2X2  AND2X2_43
timestamp 1696145522
transform 1 0 1004 0 1 2505
box -2 -3 34 103
use INVX2  INVX2_71
timestamp 1696145522
transform -1 0 1052 0 1 2505
box -2 -3 18 103
use NAND2X1  NAND2X1_133
timestamp 1696145522
transform 1 0 1052 0 1 2505
box -2 -3 26 103
use AND2X2  AND2X2_50
timestamp 1696145522
transform 1 0 1076 0 1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_294
timestamp 1696145522
transform 1 0 1108 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_635
timestamp 1696145522
transform 1 0 1140 0 1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_424
timestamp 1696145522
transform 1 0 1172 0 1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_674
timestamp 1696145522
transform -1 0 1228 0 1 2505
box -2 -3 34 103
use INVX2  INVX2_60
timestamp 1696145522
transform 1 0 1228 0 1 2505
box -2 -3 18 103
use INVX2  INVX2_44
timestamp 1696145522
transform 1 0 1244 0 1 2505
box -2 -3 18 103
use NAND2X1  NAND2X1_126
timestamp 1696145522
transform 1 0 1260 0 1 2505
box -2 -3 26 103
use BUFX4  BUFX4_149
timestamp 1696145522
transform -1 0 1316 0 1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_374
timestamp 1696145522
transform 1 0 1316 0 1 2505
box -2 -3 26 103
use BUFX4  BUFX4_153
timestamp 1696145522
transform -1 0 1372 0 1 2505
box -2 -3 34 103
use INVX8  INVX8_16
timestamp 1696145522
transform -1 0 1412 0 1 2505
box -2 -3 42 103
use NOR2X1  NOR2X1_201
timestamp 1696145522
transform 1 0 1412 0 1 2505
box -2 -3 26 103
use INVX2  INVX2_72
timestamp 1696145522
transform 1 0 1436 0 1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_410
timestamp 1696145522
transform 1 0 1452 0 1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_555
timestamp 1696145522
transform -1 0 1508 0 1 2505
box -2 -3 26 103
use FILL  FILL_25_2_0
timestamp 1696145522
transform 1 0 1508 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_2_1
timestamp 1696145522
transform 1 0 1516 0 1 2505
box -2 -3 10 103
use NOR2X1  NOR2X1_202
timestamp 1696145522
transform 1 0 1524 0 1 2505
box -2 -3 26 103
use AOI22X1  AOI22X1_11
timestamp 1696145522
transform 1 0 1548 0 1 2505
box -2 -3 42 103
use OAI21X1  OAI21X1_407
timestamp 1696145522
transform -1 0 1620 0 1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_138
timestamp 1696145522
transform -1 0 1652 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_408
timestamp 1696145522
transform 1 0 1652 0 1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_218
timestamp 1696145522
transform 1 0 1684 0 1 2505
box -2 -3 26 103
use AOI21X1  AOI21X1_293
timestamp 1696145522
transform -1 0 1740 0 1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_400
timestamp 1696145522
transform 1 0 1740 0 1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_399
timestamp 1696145522
transform -1 0 1788 0 1 2505
box -2 -3 26 103
use INVX8  INVX8_11
timestamp 1696145522
transform -1 0 1828 0 1 2505
box -2 -3 42 103
use OAI21X1  OAI21X1_409
timestamp 1696145522
transform 1 0 1828 0 1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_132
timestamp 1696145522
transform 1 0 1860 0 1 2505
box -2 -3 34 103
use BUFX4  BUFX4_144
timestamp 1696145522
transform 1 0 1892 0 1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_178
timestamp 1696145522
transform -1 0 1956 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_500
timestamp 1696145522
transform -1 0 1988 0 1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_436
timestamp 1696145522
transform 1 0 1988 0 1 2505
box -2 -3 26 103
use NOR2X1  NOR2X1_412
timestamp 1696145522
transform -1 0 2036 0 1 2505
box -2 -3 26 103
use FILL  FILL_25_3_0
timestamp 1696145522
transform -1 0 2044 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_3_1
timestamp 1696145522
transform -1 0 2052 0 1 2505
box -2 -3 10 103
use INVX1  INVX1_158
timestamp 1696145522
transform -1 0 2068 0 1 2505
box -2 -3 18 103
use AND2X2  AND2X2_27
timestamp 1696145522
transform -1 0 2100 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_362
timestamp 1696145522
transform -1 0 2132 0 1 2505
box -2 -3 34 103
use INVX1  INVX1_157
timestamp 1696145522
transform -1 0 2148 0 1 2505
box -2 -3 18 103
use NAND2X1  NAND2X1_437
timestamp 1696145522
transform 1 0 2148 0 1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_364
timestamp 1696145522
transform 1 0 2172 0 1 2505
box -2 -3 26 103
use INVX1  INVX1_126
timestamp 1696145522
transform -1 0 2212 0 1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_288
timestamp 1696145522
transform -1 0 2244 0 1 2505
box -2 -3 34 103
use INVX1  INVX1_127
timestamp 1696145522
transform -1 0 2260 0 1 2505
box -2 -3 18 103
use BUFX4  BUFX4_147
timestamp 1696145522
transform 1 0 2260 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_289
timestamp 1696145522
transform 1 0 2292 0 1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_85
timestamp 1696145522
transform -1 0 2356 0 1 2505
box -2 -3 34 103
use INVX2  INVX2_61
timestamp 1696145522
transform 1 0 2356 0 1 2505
box -2 -3 18 103
use INVX1  INVX1_198
timestamp 1696145522
transform 1 0 2372 0 1 2505
box -2 -3 18 103
use NOR2X1  NOR2X1_346
timestamp 1696145522
transform 1 0 2388 0 1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_666
timestamp 1696145522
transform -1 0 2444 0 1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_550
timestamp 1696145522
transform -1 0 2468 0 1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_236
timestamp 1696145522
transform 1 0 2468 0 1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_287
timestamp 1696145522
transform -1 0 2524 0 1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_158
timestamp 1696145522
transform -1 0 2548 0 1 2505
box -2 -3 26 103
use FILL  FILL_25_4_0
timestamp 1696145522
transform -1 0 2556 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_4_1
timestamp 1696145522
transform -1 0 2564 0 1 2505
box -2 -3 10 103
use OAI21X1  OAI21X1_243
timestamp 1696145522
transform -1 0 2596 0 1 2505
box -2 -3 34 103
use NAND3X1  NAND3X1_11
timestamp 1696145522
transform 1 0 2596 0 1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_190
timestamp 1696145522
transform 1 0 2628 0 1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_270
timestamp 1696145522
transform -1 0 2684 0 1 2505
box -2 -3 34 103
use INVX1  INVX1_108
timestamp 1696145522
transform 1 0 2684 0 1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_240
timestamp 1696145522
transform -1 0 2732 0 1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_268
timestamp 1696145522
transform -1 0 2756 0 1 2505
box -2 -3 26 103
use INVX1  INVX1_78
timestamp 1696145522
transform 1 0 2756 0 1 2505
box -2 -3 18 103
use NOR2X1  NOR2X1_111
timestamp 1696145522
transform -1 0 2796 0 1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_155
timestamp 1696145522
transform -1 0 2828 0 1 2505
box -2 -3 34 103
use INVX1  INVX1_77
timestamp 1696145522
transform -1 0 2844 0 1 2505
box -2 -3 18 103
use INVX2  INVX2_50
timestamp 1696145522
transform 1 0 2844 0 1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_147
timestamp 1696145522
transform 1 0 2860 0 1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_510
timestamp 1696145522
transform -1 0 2916 0 1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_949
timestamp 1696145522
transform -1 0 2948 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_948
timestamp 1696145522
transform 1 0 2948 0 1 2505
box -2 -3 34 103
use OAI21X1  OAI21X1_947
timestamp 1696145522
transform -1 0 3012 0 1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_46
timestamp 1696145522
transform 1 0 3012 0 1 2505
box -2 -3 34 103
use FILL  FILL_25_5_0
timestamp 1696145522
transform -1 0 3052 0 1 2505
box -2 -3 10 103
use FILL  FILL_25_5_1
timestamp 1696145522
transform -1 0 3060 0 1 2505
box -2 -3 10 103
use AND2X2  AND2X2_9
timestamp 1696145522
transform -1 0 3092 0 1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_197
timestamp 1696145522
transform -1 0 3116 0 1 2505
box -2 -3 26 103
use OAI21X1  OAI21X1_654
timestamp 1696145522
transform -1 0 3148 0 1 2505
box -2 -3 34 103
use AOI21X1  AOI21X1_284
timestamp 1696145522
transform 1 0 3148 0 1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_414
timestamp 1696145522
transform 1 0 3180 0 1 2505
box -2 -3 26 103
use NAND2X1  NAND2X1_84
timestamp 1696145522
transform 1 0 3204 0 1 2505
box -2 -3 26 103
use INVX1  INVX1_34
timestamp 1696145522
transform 1 0 3228 0 1 2505
box -2 -3 18 103
use AOI21X1  AOI21X1_413
timestamp 1696145522
transform -1 0 3276 0 1 2505
box -2 -3 34 103
use NOR2X1  NOR2X1_2
timestamp 1696145522
transform -1 0 3300 0 1 2505
box -2 -3 26 103
use INVX1  INVX1_1
timestamp 1696145522
transform -1 0 3316 0 1 2505
box -2 -3 18 103
use OAI21X1  OAI21X1_25
timestamp 1696145522
transform 1 0 3316 0 1 2505
box -2 -3 34 103
use NAND2X1  NAND2X1_3
timestamp 1696145522
transform 1 0 3348 0 1 2505
box -2 -3 26 103
use XNOR2X1  XNOR2X1_3
timestamp 1696145522
transform -1 0 3428 0 1 2505
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_27
timestamp 1696145522
transform 1 0 3428 0 1 2505
box -2 -3 98 103
use BUFX2  BUFX2_29
timestamp 1696145522
transform 1 0 3524 0 1 2505
box -2 -3 26 103
use FILL  FILL_26_1
timestamp 1696145522
transform 1 0 3548 0 1 2505
box -2 -3 10 103
use FILL  FILL_26_2
timestamp 1696145522
transform 1 0 3556 0 1 2505
box -2 -3 10 103
use INVX1  INVX1_235
timestamp 1696145522
transform 1 0 4 0 -1 2705
box -2 -3 18 103
use OAI22X1  OAI22X1_25
timestamp 1696145522
transform -1 0 60 0 -1 2705
box -2 -3 42 103
use NOR2X1  NOR2X1_318
timestamp 1696145522
transform 1 0 60 0 -1 2705
box -2 -3 26 103
use INVX1  INVX1_230
timestamp 1696145522
transform -1 0 100 0 -1 2705
box -2 -3 18 103
use NOR2X1  NOR2X1_319
timestamp 1696145522
transform 1 0 100 0 -1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_579
timestamp 1696145522
transform 1 0 124 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_574
timestamp 1696145522
transform 1 0 156 0 -1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_320
timestamp 1696145522
transform 1 0 188 0 -1 2705
box -2 -3 26 103
use NOR2X1  NOR2X1_322
timestamp 1696145522
transform 1 0 212 0 -1 2705
box -2 -3 26 103
use NOR2X1  NOR2X1_305
timestamp 1696145522
transform -1 0 260 0 -1 2705
box -2 -3 26 103
use AOI21X1  AOI21X1_232
timestamp 1696145522
transform 1 0 260 0 -1 2705
box -2 -3 34 103
use AOI22X1  AOI22X1_25
timestamp 1696145522
transform 1 0 292 0 -1 2705
box -2 -3 42 103
use NOR2X1  NOR2X1_304
timestamp 1696145522
transform -1 0 356 0 -1 2705
box -2 -3 26 103
use NOR2X1  NOR2X1_306
timestamp 1696145522
transform 1 0 356 0 -1 2705
box -2 -3 26 103
use AOI22X1  AOI22X1_24
timestamp 1696145522
transform -1 0 420 0 -1 2705
box -2 -3 42 103
use NAND2X1  NAND2X1_516
timestamp 1696145522
transform 1 0 420 0 -1 2705
box -2 -3 26 103
use NOR2X1  NOR2X1_356
timestamp 1696145522
transform 1 0 444 0 -1 2705
box -2 -3 26 103
use INVX4  INVX4_24
timestamp 1696145522
transform 1 0 468 0 -1 2705
box -2 -3 26 103
use FILL  FILL_26_0_0
timestamp 1696145522
transform 1 0 492 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_0_1
timestamp 1696145522
transform 1 0 500 0 -1 2705
box -2 -3 10 103
use INVX1  INVX1_251
timestamp 1696145522
transform 1 0 508 0 -1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_611
timestamp 1696145522
transform 1 0 524 0 -1 2705
box -2 -3 34 103
use OAI22X1  OAI22X1_20
timestamp 1696145522
transform 1 0 556 0 -1 2705
box -2 -3 42 103
use INVX2  INVX2_53
timestamp 1696145522
transform -1 0 612 0 -1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_609
timestamp 1696145522
transform -1 0 644 0 -1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_262
timestamp 1696145522
transform 1 0 644 0 -1 2705
box -2 -3 34 103
use INVX1  INVX1_260
timestamp 1696145522
transform 1 0 676 0 -1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_623
timestamp 1696145522
transform 1 0 692 0 -1 2705
box -2 -3 34 103
use OR2X2  OR2X2_38
timestamp 1696145522
transform 1 0 724 0 -1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_411
timestamp 1696145522
transform 1 0 756 0 -1 2705
box -2 -3 26 103
use NOR2X1  NOR2X1_367
timestamp 1696145522
transform -1 0 804 0 -1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_521
timestamp 1696145522
transform -1 0 828 0 -1 2705
box -2 -3 26 103
use INVX1  INVX1_259
timestamp 1696145522
transform 1 0 828 0 -1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_620
timestamp 1696145522
transform 1 0 844 0 -1 2705
box -2 -3 34 103
use INVX2  INVX2_91
timestamp 1696145522
transform 1 0 876 0 -1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_626
timestamp 1696145522
transform 1 0 892 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_627
timestamp 1696145522
transform -1 0 956 0 -1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_267
timestamp 1696145522
transform 1 0 956 0 -1 2705
box -2 -3 34 103
use FILL  FILL_26_1_0
timestamp 1696145522
transform 1 0 988 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_1_1
timestamp 1696145522
transform 1 0 996 0 -1 2705
box -2 -3 10 103
use AOI21X1  AOI21X1_271
timestamp 1696145522
transform 1 0 1004 0 -1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_525
timestamp 1696145522
transform -1 0 1060 0 -1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_537
timestamp 1696145522
transform -1 0 1084 0 -1 2705
box -2 -3 26 103
use AOI21X1  AOI21X1_273
timestamp 1696145522
transform 1 0 1084 0 -1 2705
box -2 -3 34 103
use NAND3X1  NAND3X1_33
timestamp 1696145522
transform 1 0 1116 0 -1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_275
timestamp 1696145522
transform 1 0 1148 0 -1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_528
timestamp 1696145522
transform -1 0 1204 0 -1 2705
box -2 -3 26 103
use NOR2X1  NOR2X1_371
timestamp 1696145522
transform -1 0 1228 0 -1 2705
box -2 -3 26 103
use INVX2  INVX2_42
timestamp 1696145522
transform -1 0 1244 0 -1 2705
box -2 -3 18 103
use AND2X2  AND2X2_44
timestamp 1696145522
transform -1 0 1276 0 -1 2705
box -2 -3 34 103
use BUFX4  BUFX4_145
timestamp 1696145522
transform -1 0 1308 0 -1 2705
box -2 -3 34 103
use INVX2  INVX2_54
timestamp 1696145522
transform -1 0 1324 0 -1 2705
box -2 -3 18 103
use BUFX4  BUFX4_56
timestamp 1696145522
transform -1 0 1356 0 -1 2705
box -2 -3 34 103
use NAND3X1  NAND3X1_30
timestamp 1696145522
transform 1 0 1356 0 -1 2705
box -2 -3 34 103
use BUFX4  BUFX4_64
timestamp 1696145522
transform -1 0 1420 0 -1 2705
box -2 -3 34 103
use BUFX4  BUFX4_146
timestamp 1696145522
transform 1 0 1420 0 -1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_553
timestamp 1696145522
transform -1 0 1476 0 -1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_672
timestamp 1696145522
transform -1 0 1508 0 -1 2705
box -2 -3 34 103
use FILL  FILL_26_2_0
timestamp 1696145522
transform 1 0 1508 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_2_1
timestamp 1696145522
transform 1 0 1516 0 -1 2705
box -2 -3 10 103
use NOR2X1  NOR2X1_189
timestamp 1696145522
transform 1 0 1524 0 -1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_389
timestamp 1696145522
transform 1 0 1548 0 -1 2705
box -2 -3 34 103
use AOI22X1  AOI22X1_10
timestamp 1696145522
transform -1 0 1620 0 -1 2705
box -2 -3 42 103
use NAND2X1  NAND2X1_554
timestamp 1696145522
transform -1 0 1644 0 -1 2705
box -2 -3 26 103
use AOI21X1  AOI21X1_125
timestamp 1696145522
transform -1 0 1676 0 -1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_179
timestamp 1696145522
transform -1 0 1700 0 -1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_389
timestamp 1696145522
transform 1 0 1700 0 -1 2705
box -2 -3 26 103
use NOR2X1  NOR2X1_185
timestamp 1696145522
transform 1 0 1724 0 -1 2705
box -2 -3 26 103
use AOI21X1  AOI21X1_117
timestamp 1696145522
transform -1 0 1780 0 -1 2705
box -2 -3 34 103
use AND2X2  AND2X2_19
timestamp 1696145522
transform 1 0 1780 0 -1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_130
timestamp 1696145522
transform 1 0 1812 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_392
timestamp 1696145522
transform -1 0 1876 0 -1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_382
timestamp 1696145522
transform -1 0 1900 0 -1 2705
box -2 -3 26 103
use NOR2X1  NOR2X1_191
timestamp 1696145522
transform -1 0 1924 0 -1 2705
box -2 -3 26 103
use AND2X2  AND2X2_17
timestamp 1696145522
transform -1 0 1956 0 -1 2705
box -2 -3 34 103
use INVX1  INVX1_163
timestamp 1696145522
transform -1 0 1972 0 -1 2705
box -2 -3 18 103
use BUFX4  BUFX4_61
timestamp 1696145522
transform -1 0 2004 0 -1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_282
timestamp 1696145522
transform 1 0 2004 0 -1 2705
box -2 -3 26 103
use FILL  FILL_26_3_0
timestamp 1696145522
transform -1 0 2036 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_3_1
timestamp 1696145522
transform -1 0 2044 0 -1 2705
box -2 -3 10 103
use NAND2X1  NAND2X1_469
timestamp 1696145522
transform -1 0 2068 0 -1 2705
box -2 -3 26 103
use INVX1  INVX1_154
timestamp 1696145522
transform 1 0 2068 0 -1 2705
box -2 -3 18 103
use AOI21X1  AOI21X1_112
timestamp 1696145522
transform 1 0 2084 0 -1 2705
box -2 -3 34 103
use INVX1  INVX1_155
timestamp 1696145522
transform -1 0 2132 0 -1 2705
box -2 -3 18 103
use AOI21X1  AOI21X1_118
timestamp 1696145522
transform -1 0 2164 0 -1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_362
timestamp 1696145522
transform 1 0 2164 0 -1 2705
box -2 -3 26 103
use AOI21X1  AOI21X1_115
timestamp 1696145522
transform 1 0 2188 0 -1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_137
timestamp 1696145522
transform 1 0 2220 0 -1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_184
timestamp 1696145522
transform 1 0 2252 0 -1 2705
box -2 -3 26 103
use NOR2X1  NOR2X1_183
timestamp 1696145522
transform 1 0 2276 0 -1 2705
box -2 -3 26 103
use NOR2X1  NOR2X1_182
timestamp 1696145522
transform 1 0 2300 0 -1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_667
timestamp 1696145522
transform -1 0 2356 0 -1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_421
timestamp 1696145522
transform 1 0 2356 0 -1 2705
box -2 -3 26 103
use NOR2X1  NOR2X1_420
timestamp 1696145522
transform 1 0 2380 0 -1 2705
box -2 -3 26 103
use AND2X2  AND2X2_15
timestamp 1696145522
transform 1 0 2404 0 -1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_165
timestamp 1696145522
transform -1 0 2468 0 -1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_435
timestamp 1696145522
transform -1 0 2492 0 -1 2705
box -2 -3 26 103
use INVX1  INVX1_153
timestamp 1696145522
transform 1 0 2492 0 -1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_359
timestamp 1696145522
transform -1 0 2540 0 -1 2705
box -2 -3 34 103
use FILL  FILL_26_4_0
timestamp 1696145522
transform 1 0 2540 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_4_1
timestamp 1696145522
transform 1 0 2548 0 -1 2705
box -2 -3 10 103
use NOR2X1  NOR2X1_245
timestamp 1696145522
transform 1 0 2556 0 -1 2705
box -2 -3 26 103
use OR2X2  OR2X2_17
timestamp 1696145522
transform -1 0 2612 0 -1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_291
timestamp 1696145522
transform 1 0 2612 0 -1 2705
box -2 -3 34 103
use INVX1  INVX1_283
timestamp 1696145522
transform -1 0 2660 0 -1 2705
box -2 -3 18 103
use NAND2X1  NAND2X1_307
timestamp 1696145522
transform 1 0 2660 0 -1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_665
timestamp 1696145522
transform -1 0 2716 0 -1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_548
timestamp 1696145522
transform -1 0 2740 0 -1 2705
box -2 -3 26 103
use AOI21X1  AOI21X1_80
timestamp 1696145522
transform 1 0 2740 0 -1 2705
box -2 -3 34 103
use OAI22X1  OAI22X1_3
timestamp 1696145522
transform 1 0 2772 0 -1 2705
box -2 -3 42 103
use AOI21X1  AOI21X1_82
timestamp 1696145522
transform 1 0 2812 0 -1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_155
timestamp 1696145522
transform -1 0 2868 0 -1 2705
box -2 -3 26 103
use AOI22X1  AOI22X1_6
timestamp 1696145522
transform 1 0 2868 0 -1 2705
box -2 -3 42 103
use NAND2X1  NAND2X1_289
timestamp 1696145522
transform -1 0 2932 0 -1 2705
box -2 -3 26 103
use AOI21X1  AOI21X1_65
timestamp 1696145522
transform 1 0 2932 0 -1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_69
timestamp 1696145522
transform 1 0 2964 0 -1 2705
box -2 -3 34 103
use AOI22X1  AOI22X1_3
timestamp 1696145522
transform -1 0 3036 0 -1 2705
box -2 -3 42 103
use FILL  FILL_26_5_0
timestamp 1696145522
transform -1 0 3044 0 -1 2705
box -2 -3 10 103
use FILL  FILL_26_5_1
timestamp 1696145522
transform -1 0 3052 0 -1 2705
box -2 -3 10 103
use AND2X2  AND2X2_4
timestamp 1696145522
transform -1 0 3084 0 -1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_92
timestamp 1696145522
transform -1 0 3116 0 -1 2705
box -2 -3 34 103
use INVX2  INVX2_35
timestamp 1696145522
transform 1 0 3116 0 -1 2705
box -2 -3 18 103
use NAND2X1  NAND2X1_193
timestamp 1696145522
transform -1 0 3156 0 -1 2705
box -2 -3 26 103
use NOR2X1  NOR2X1_95
timestamp 1696145522
transform -1 0 3180 0 -1 2705
box -2 -3 26 103
use NOR2X1  NOR2X1_105
timestamp 1696145522
transform -1 0 3204 0 -1 2705
box -2 -3 26 103
use NOR2X1  NOR2X1_3
timestamp 1696145522
transform 1 0 3204 0 -1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_204
timestamp 1696145522
transform -1 0 3252 0 -1 2705
box -2 -3 26 103
use AOI21X1  AOI21X1_34
timestamp 1696145522
transform 1 0 3252 0 -1 2705
box -2 -3 34 103
use XNOR2X1  XNOR2X1_2
timestamp 1696145522
transform 1 0 3284 0 -1 2705
box -2 -3 58 103
use AOI21X1  AOI21X1_1
timestamp 1696145522
transform 1 0 3340 0 -1 2705
box -2 -3 34 103
use INVX1  INVX1_329
timestamp 1696145522
transform -1 0 3388 0 -1 2705
box -2 -3 18 103
use NAND2X1  NAND2X1_2
timestamp 1696145522
transform -1 0 3412 0 -1 2705
box -2 -3 26 103
use NOR2X1  NOR2X1_1
timestamp 1696145522
transform -1 0 3436 0 -1 2705
box -2 -3 26 103
use INVX1  INVX1_326
timestamp 1696145522
transform 1 0 3436 0 -1 2705
box -2 -3 18 103
use NAND2X1  NAND2X1_1
timestamp 1696145522
transform 1 0 3452 0 -1 2705
box -2 -3 26 103
use INVX2  INVX2_1
timestamp 1696145522
transform -1 0 3492 0 -1 2705
box -2 -3 18 103
use XNOR2X1  XNOR2X1_1
timestamp 1696145522
transform -1 0 3548 0 -1 2705
box -2 -3 58 103
use FILL  FILL_27_1
timestamp 1696145522
transform -1 0 3556 0 -1 2705
box -2 -3 10 103
use FILL  FILL_27_2
timestamp 1696145522
transform -1 0 3564 0 -1 2705
box -2 -3 10 103
use INVX2  INVX2_85
timestamp 1696145522
transform 1 0 4 0 1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_657
timestamp 1696145522
transform 1 0 20 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_584
timestamp 1696145522
transform 1 0 52 0 1 2705
box -2 -3 34 103
use INVX1  INVX1_240
timestamp 1696145522
transform 1 0 84 0 1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_585
timestamp 1696145522
transform -1 0 132 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_575
timestamp 1696145522
transform 1 0 132 0 1 2705
box -2 -3 34 103
use INVX1  INVX1_237
timestamp 1696145522
transform -1 0 180 0 1 2705
box -2 -3 18 103
use NAND2X1  NAND2X1_512
timestamp 1696145522
transform 1 0 180 0 1 2705
box -2 -3 26 103
use NOR2X1  NOR2X1_324
timestamp 1696145522
transform -1 0 228 0 1 2705
box -2 -3 26 103
use NOR2X1  NOR2X1_323
timestamp 1696145522
transform 1 0 228 0 1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_573
timestamp 1696145522
transform -1 0 284 0 1 2705
box -2 -3 34 103
use INVX2  INVX2_82
timestamp 1696145522
transform -1 0 300 0 1 2705
box -2 -3 18 103
use AOI21X1  AOI21X1_230
timestamp 1696145522
transform 1 0 300 0 1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_325
timestamp 1696145522
transform -1 0 356 0 1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_610
timestamp 1696145522
transform 1 0 356 0 1 2705
box -2 -3 34 103
use INVX1  INVX1_253
timestamp 1696145522
transform -1 0 404 0 1 2705
box -2 -3 18 103
use INVX2  INVX2_81
timestamp 1696145522
transform -1 0 420 0 1 2705
box -2 -3 18 103
use AOI21X1  AOI21X1_259
timestamp 1696145522
transform -1 0 452 0 1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_266
timestamp 1696145522
transform 1 0 452 0 1 2705
box -2 -3 34 103
use FILL  FILL_27_0_0
timestamp 1696145522
transform -1 0 492 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_0_1
timestamp 1696145522
transform -1 0 500 0 1 2705
box -2 -3 10 103
use INVX2  INVX2_89
timestamp 1696145522
transform -1 0 516 0 1 2705
box -2 -3 18 103
use INVX1  INVX1_257
timestamp 1696145522
transform -1 0 532 0 1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_619
timestamp 1696145522
transform -1 0 564 0 1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_366
timestamp 1696145522
transform -1 0 588 0 1 2705
box -2 -3 26 103
use INVX2  INVX2_88
timestamp 1696145522
transform -1 0 604 0 1 2705
box -2 -3 18 103
use INVX2  INVX2_80
timestamp 1696145522
transform 1 0 604 0 1 2705
box -2 -3 18 103
use AOI21X1  AOI21X1_251
timestamp 1696145522
transform -1 0 652 0 1 2705
box -2 -3 34 103
use INVX1  INVX1_248
timestamp 1696145522
transform -1 0 668 0 1 2705
box -2 -3 18 103
use AOI21X1  AOI21X1_264
timestamp 1696145522
transform 1 0 668 0 1 2705
box -2 -3 34 103
use INVX1  INVX1_258
timestamp 1696145522
transform 1 0 700 0 1 2705
box -2 -3 18 103
use AOI21X1  AOI21X1_265
timestamp 1696145522
transform 1 0 716 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_621
timestamp 1696145522
transform 1 0 748 0 1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_219
timestamp 1696145522
transform 1 0 780 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_566
timestamp 1696145522
transform 1 0 812 0 1 2705
box -2 -3 34 103
use OAI22X1  OAI22X1_22
timestamp 1696145522
transform -1 0 884 0 1 2705
box -2 -3 42 103
use AOI21X1  AOI21X1_269
timestamp 1696145522
transform -1 0 916 0 1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_205
timestamp 1696145522
transform -1 0 948 0 1 2705
box -2 -3 34 103
use NAND3X1  NAND3X1_38
timestamp 1696145522
transform 1 0 948 0 1 2705
box -2 -3 34 103
use NAND3X1  NAND3X1_37
timestamp 1696145522
transform -1 0 1012 0 1 2705
box -2 -3 34 103
use FILL  FILL_27_1_0
timestamp 1696145522
transform 1 0 1012 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_1_1
timestamp 1696145522
transform 1 0 1020 0 1 2705
box -2 -3 10 103
use INVX1  INVX1_236
timestamp 1696145522
transform 1 0 1028 0 1 2705
box -2 -3 18 103
use AOI21X1  AOI21X1_225
timestamp 1696145522
transform -1 0 1076 0 1 2705
box -2 -3 34 103
use NAND3X1  NAND3X1_39
timestamp 1696145522
transform -1 0 1108 0 1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_484
timestamp 1696145522
transform 1 0 1108 0 1 2705
box -2 -3 26 103
use INVX2  INVX2_41
timestamp 1696145522
transform -1 0 1148 0 1 2705
box -2 -3 18 103
use AOI21X1  AOI21X1_276
timestamp 1696145522
transform 1 0 1148 0 1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_270
timestamp 1696145522
transform 1 0 1180 0 1 2705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_64
timestamp 1696145522
transform 1 0 1204 0 1 2705
box -2 -3 98 103
use NOR2X1  NOR2X1_375
timestamp 1696145522
transform -1 0 1324 0 1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_458
timestamp 1696145522
transform -1 0 1348 0 1 2705
box -2 -3 26 103
use AOI22X1  AOI22X1_21
timestamp 1696145522
transform 1 0 1348 0 1 2705
box -2 -3 42 103
use INVX2  INVX2_52
timestamp 1696145522
transform -1 0 1404 0 1 2705
box -2 -3 18 103
use NOR2X1  NOR2X1_370
timestamp 1696145522
transform -1 0 1428 0 1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_634
timestamp 1696145522
transform -1 0 1460 0 1 2705
box -2 -3 34 103
use AND2X2  AND2X2_38
timestamp 1696145522
transform 1 0 1460 0 1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_188
timestamp 1696145522
transform 1 0 1492 0 1 2705
box -2 -3 26 103
use FILL  FILL_27_2_0
timestamp 1696145522
transform 1 0 1516 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_2_1
timestamp 1696145522
transform 1 0 1524 0 1 2705
box -2 -3 10 103
use INVX1  INVX1_161
timestamp 1696145522
transform 1 0 1532 0 1 2705
box -2 -3 18 103
use NOR2X1  NOR2X1_190
timestamp 1696145522
transform 1 0 1548 0 1 2705
box -2 -3 26 103
use INVX2  INVX2_55
timestamp 1696145522
transform -1 0 1588 0 1 2705
box -2 -3 18 103
use NAND2X1  NAND2X1_383
timestamp 1696145522
transform 1 0 1588 0 1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_394
timestamp 1696145522
transform -1 0 1644 0 1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_178
timestamp 1696145522
transform 1 0 1644 0 1 2705
box -2 -3 26 103
use INVX1  INVX1_152
timestamp 1696145522
transform -1 0 1684 0 1 2705
box -2 -3 18 103
use NAND2X1  NAND2X1_376
timestamp 1696145522
transform -1 0 1708 0 1 2705
box -2 -3 26 103
use NOR2X1  NOR2X1_180
timestamp 1696145522
transform -1 0 1732 0 1 2705
box -2 -3 26 103
use INVX1  INVX1_169
timestamp 1696145522
transform 1 0 1732 0 1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_395
timestamp 1696145522
transform -1 0 1780 0 1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_203
timestamp 1696145522
transform 1 0 1780 0 1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_384
timestamp 1696145522
transform 1 0 1804 0 1 2705
box -2 -3 26 103
use BUFX4  BUFX4_94
timestamp 1696145522
transform -1 0 1860 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_381
timestamp 1696145522
transform 1 0 1860 0 1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_192
timestamp 1696145522
transform 1 0 1892 0 1 2705
box -2 -3 26 103
use AND2X2  AND2X2_16
timestamp 1696145522
transform 1 0 1916 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_380
timestamp 1696145522
transform -1 0 1980 0 1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_123
timestamp 1696145522
transform 1 0 1980 0 1 2705
box -2 -3 34 103
use FILL  FILL_27_3_0
timestamp 1696145522
transform -1 0 2020 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_3_1
timestamp 1696145522
transform -1 0 2028 0 1 2705
box -2 -3 10 103
use BUFX4  BUFX4_93
timestamp 1696145522
transform -1 0 2060 0 1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_114
timestamp 1696145522
transform 1 0 2060 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_363
timestamp 1696145522
transform -1 0 2124 0 1 2705
box -2 -3 34 103
use INVX1  INVX1_156
timestamp 1696145522
transform 1 0 2124 0 1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_364
timestamp 1696145522
transform 1 0 2140 0 1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_164
timestamp 1696145522
transform 1 0 2172 0 1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_547
timestamp 1696145522
transform 1 0 2196 0 1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_664
timestamp 1696145522
transform -1 0 2252 0 1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_98
timestamp 1696145522
transform -1 0 2284 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_331
timestamp 1696145522
transform -1 0 2316 0 1 2705
box -2 -3 34 103
use INVX1  INVX1_144
timestamp 1696145522
transform -1 0 2332 0 1 2705
box -2 -3 18 103
use AOI21X1  AOI21X1_91
timestamp 1696145522
transform -1 0 2364 0 1 2705
box -2 -3 34 103
use INVX2  INVX2_65
timestamp 1696145522
transform -1 0 2380 0 1 2705
box -2 -3 18 103
use XNOR2X1  XNOR2X1_32
timestamp 1696145522
transform 1 0 2380 0 1 2705
box -2 -3 58 103
use AOI21X1  AOI21X1_95
timestamp 1696145522
transform -1 0 2468 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_472
timestamp 1696145522
transform -1 0 2500 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_358
timestamp 1696145522
transform -1 0 2532 0 1 2705
box -2 -3 34 103
use FILL  FILL_27_4_0
timestamp 1696145522
transform -1 0 2540 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_4_1
timestamp 1696145522
transform -1 0 2548 0 1 2705
box -2 -3 10 103
use OAI21X1  OAI21X1_284
timestamp 1696145522
transform -1 0 2580 0 1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_157
timestamp 1696145522
transform -1 0 2604 0 1 2705
box -2 -3 26 103
use AOI21X1  AOI21X1_84
timestamp 1696145522
transform -1 0 2636 0 1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_156
timestamp 1696145522
transform -1 0 2660 0 1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_264
timestamp 1696145522
transform 1 0 2660 0 1 2705
box -2 -3 34 103
use XNOR2X1  XNOR2X1_31
timestamp 1696145522
transform 1 0 2692 0 1 2705
box -2 -3 58 103
use AOI21X1  AOI21X1_73
timestamp 1696145522
transform 1 0 2748 0 1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_134
timestamp 1696145522
transform 1 0 2780 0 1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_286
timestamp 1696145522
transform 1 0 2804 0 1 2705
box -2 -3 34 103
use INVX2  INVX2_62
timestamp 1696145522
transform 1 0 2836 0 1 2705
box -2 -3 18 103
use NAND2X1  NAND2X1_287
timestamp 1696145522
transform 1 0 2852 0 1 2705
box -2 -3 26 103
use INVX1  INVX1_116
timestamp 1696145522
transform -1 0 2892 0 1 2705
box -2 -3 18 103
use BUFX4  BUFX4_95
timestamp 1696145522
transform 1 0 2892 0 1 2705
box -2 -3 34 103
use NAND2X1  NAND2X1_288
timestamp 1696145522
transform -1 0 2948 0 1 2705
box -2 -3 26 103
use NOR2X1  NOR2X1_130
timestamp 1696145522
transform 1 0 2948 0 1 2705
box -2 -3 26 103
use AOI22X1  AOI22X1_2
timestamp 1696145522
transform 1 0 2972 0 1 2705
box -2 -3 42 103
use NAND3X1  NAND3X1_3
timestamp 1696145522
transform -1 0 3044 0 1 2705
box -2 -3 34 103
use FILL  FILL_27_5_0
timestamp 1696145522
transform -1 0 3052 0 1 2705
box -2 -3 10 103
use FILL  FILL_27_5_1
timestamp 1696145522
transform -1 0 3060 0 1 2705
box -2 -3 10 103
use AOI21X1  AOI21X1_45
timestamp 1696145522
transform -1 0 3092 0 1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_285
timestamp 1696145522
transform -1 0 3124 0 1 2705
box -2 -3 34 103
use INVX1  INVX1_76
timestamp 1696145522
transform -1 0 3140 0 1 2705
box -2 -3 18 103
use OAI21X1  OAI21X1_150
timestamp 1696145522
transform -1 0 3172 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_149
timestamp 1696145522
transform 1 0 3172 0 1 2705
box -2 -3 34 103
use AOI21X1  AOI21X1_56
timestamp 1696145522
transform -1 0 3236 0 1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_119
timestamp 1696145522
transform 1 0 3236 0 1 2705
box -2 -3 26 103
use NAND2X1  NAND2X1_206
timestamp 1696145522
transform -1 0 3284 0 1 2705
box -2 -3 26 103
use OAI21X1  OAI21X1_173
timestamp 1696145522
transform -1 0 3316 0 1 2705
box -2 -3 34 103
use INVX1  INVX1_2
timestamp 1696145522
transform -1 0 3332 0 1 2705
box -2 -3 18 103
use AND2X2  AND2X2_5
timestamp 1696145522
transform -1 0 3364 0 1 2705
box -2 -3 34 103
use AND2X2  AND2X2_2
timestamp 1696145522
transform -1 0 3396 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_172
timestamp 1696145522
transform -1 0 3428 0 1 2705
box -2 -3 34 103
use OAI21X1  OAI21X1_937
timestamp 1696145522
transform -1 0 3460 0 1 2705
box -2 -3 34 103
use NOR2X1  NOR2X1_504
timestamp 1696145522
transform 1 0 3460 0 1 2705
box -2 -3 26 103
use NOR2X1  NOR2X1_508
timestamp 1696145522
transform 1 0 3484 0 1 2705
box -2 -3 26 103
use AND2X2  AND2X2_74
timestamp 1696145522
transform 1 0 3508 0 1 2705
box -2 -3 34 103
use BUFX2  BUFX2_67
timestamp 1696145522
transform 1 0 3540 0 1 2705
box -2 -3 26 103
use NOR2X1  NOR2X1_416
timestamp 1696145522
transform 1 0 4 0 -1 2905
box -2 -3 26 103
use INVX1  INVX1_242
timestamp 1696145522
transform 1 0 28 0 -1 2905
box -2 -3 18 103
use NOR2X1  NOR2X1_337
timestamp 1696145522
transform -1 0 68 0 -1 2905
box -2 -3 26 103
use NOR2X1  NOR2X1_349
timestamp 1696145522
transform -1 0 92 0 -1 2905
box -2 -3 26 103
use NOR2X1  NOR2X1_338
timestamp 1696145522
transform 1 0 92 0 -1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_601
timestamp 1696145522
transform -1 0 148 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_658
timestamp 1696145522
transform -1 0 180 0 -1 2905
box -2 -3 34 103
use INVX1  INVX1_249
timestamp 1696145522
transform -1 0 196 0 -1 2905
box -2 -3 18 103
use INVX1  INVX1_243
timestamp 1696145522
transform 1 0 196 0 -1 2905
box -2 -3 18 103
use NOR2X1  NOR2X1_345
timestamp 1696145522
transform -1 0 236 0 -1 2905
box -2 -3 26 103
use INVX1  INVX1_241
timestamp 1696145522
transform 1 0 236 0 -1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_596
timestamp 1696145522
transform 1 0 252 0 -1 2905
box -2 -3 34 103
use INVX1  INVX1_246
timestamp 1696145522
transform 1 0 284 0 -1 2905
box -2 -3 18 103
use AOI21X1  AOI21X1_247
timestamp 1696145522
transform -1 0 332 0 -1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_511
timestamp 1696145522
transform 1 0 332 0 -1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_594
timestamp 1696145522
transform -1 0 388 0 -1 2905
box -2 -3 34 103
use OAI22X1  OAI22X1_17
timestamp 1696145522
transform 1 0 388 0 -1 2905
box -2 -3 42 103
use NOR2X1  NOR2X1_333
timestamp 1696145522
transform 1 0 428 0 -1 2905
box -2 -3 26 103
use NOR2X1  NOR2X1_334
timestamp 1696145522
transform -1 0 476 0 -1 2905
box -2 -3 26 103
use FILL  FILL_28_0_0
timestamp 1696145522
transform -1 0 484 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_0_1
timestamp 1696145522
transform -1 0 492 0 -1 2905
box -2 -3 10 103
use OAI21X1  OAI21X1_663
timestamp 1696145522
transform -1 0 524 0 -1 2905
box -2 -3 34 103
use AND2X2  AND2X2_49
timestamp 1696145522
transform -1 0 556 0 -1 2905
box -2 -3 34 103
use AOI21X1  AOI21X1_249
timestamp 1696145522
transform -1 0 588 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_600
timestamp 1696145522
transform -1 0 620 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_597
timestamp 1696145522
transform -1 0 652 0 -1 2905
box -2 -3 34 103
use INVX1  INVX1_247
timestamp 1696145522
transform 1 0 652 0 -1 2905
box -2 -3 18 103
use NAND2X1  NAND2X1_491
timestamp 1696145522
transform 1 0 668 0 -1 2905
box -2 -3 26 103
use NOR2X1  NOR2X1_313
timestamp 1696145522
transform 1 0 692 0 -1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_543
timestamp 1696145522
transform -1 0 740 0 -1 2905
box -2 -3 26 103
use AOI21X1  AOI21X1_218
timestamp 1696145522
transform -1 0 772 0 -1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_298
timestamp 1696145522
transform -1 0 796 0 -1 2905
box -2 -3 26 103
use INVX2  INVX2_40
timestamp 1696145522
transform -1 0 812 0 -1 2905
box -2 -3 18 103
use NOR2X1  NOR2X1_290
timestamp 1696145522
transform -1 0 836 0 -1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_542
timestamp 1696145522
transform -1 0 868 0 -1 2905
box -2 -3 34 103
use OAI22X1  OAI22X1_13
timestamp 1696145522
transform -1 0 908 0 -1 2905
box -2 -3 42 103
use OAI21X1  OAI21X1_599
timestamp 1696145522
transform -1 0 940 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_565
timestamp 1696145522
transform -1 0 972 0 -1 2905
box -2 -3 34 103
use INVX1  INVX1_233
timestamp 1696145522
transform -1 0 988 0 -1 2905
box -2 -3 18 103
use FILL  FILL_28_1_0
timestamp 1696145522
transform 1 0 988 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_1_1
timestamp 1696145522
transform 1 0 996 0 -1 2905
box -2 -3 10 103
use AOI21X1  AOI21X1_272
timestamp 1696145522
transform 1 0 1004 0 -1 2905
box -2 -3 34 103
use AOI21X1  AOI21X1_217
timestamp 1696145522
transform -1 0 1068 0 -1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_369
timestamp 1696145522
transform 1 0 1068 0 -1 2905
box -2 -3 26 103
use INVX1  INVX1_231
timestamp 1696145522
transform -1 0 1108 0 -1 2905
box -2 -3 18 103
use OAI22X1  OAI22X1_11
timestamp 1696145522
transform -1 0 1148 0 -1 2905
box -2 -3 42 103
use NOR2X1  NOR2X1_262
timestamp 1696145522
transform 1 0 1148 0 -1 2905
box -2 -3 26 103
use OAI22X1  OAI22X1_26
timestamp 1696145522
transform 1 0 1172 0 -1 2905
box -2 -3 42 103
use NAND2X1  NAND2X1_461
timestamp 1696145522
transform -1 0 1236 0 -1 2905
box -2 -3 26 103
use INVX2  INVX2_77
timestamp 1696145522
transform -1 0 1252 0 -1 2905
box -2 -3 18 103
use NOR2X1  NOR2X1_271
timestamp 1696145522
transform 1 0 1252 0 -1 2905
box -2 -3 26 103
use INVX1  INVX1_214
timestamp 1696145522
transform 1 0 1276 0 -1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_517
timestamp 1696145522
transform -1 0 1324 0 -1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_541
timestamp 1696145522
transform 1 0 1324 0 -1 2905
box -2 -3 26 103
use NOR2X1  NOR2X1_256
timestamp 1696145522
transform 1 0 1348 0 -1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_495
timestamp 1696145522
transform 1 0 1372 0 -1 2905
box -2 -3 34 103
use AOI21X1  AOI21X1_179
timestamp 1696145522
transform -1 0 1436 0 -1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_265
timestamp 1696145522
transform -1 0 1460 0 -1 2905
box -2 -3 26 103
use AOI22X1  AOI22X1_20
timestamp 1696145522
transform 1 0 1460 0 -1 2905
box -2 -3 42 103
use FILL  FILL_28_2_0
timestamp 1696145522
transform 1 0 1500 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_2_1
timestamp 1696145522
transform 1 0 1508 0 -1 2905
box -2 -3 10 103
use AND2X2  AND2X2_29
timestamp 1696145522
transform 1 0 1516 0 -1 2905
box -2 -3 34 103
use AOI21X1  AOI21X1_248
timestamp 1696145522
transform -1 0 1580 0 -1 2905
box -2 -3 34 103
use XNOR2X1  XNOR2X1_36
timestamp 1696145522
transform 1 0 1580 0 -1 2905
box -2 -3 58 103
use AOI22X1  AOI22X1_18
timestamp 1696145522
transform 1 0 1636 0 -1 2905
box -2 -3 42 103
use INVX1  INVX1_202
timestamp 1696145522
transform -1 0 1692 0 -1 2905
box -2 -3 18 103
use INVX2  INVX2_69
timestamp 1696145522
transform -1 0 1708 0 -1 2905
box -2 -3 18 103
use AOI21X1  AOI21X1_126
timestamp 1696145522
transform -1 0 1740 0 -1 2905
box -2 -3 34 103
use INVX1  INVX1_201
timestamp 1696145522
transform 1 0 1740 0 -1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_393
timestamp 1696145522
transform -1 0 1788 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_486
timestamp 1696145522
transform -1 0 1820 0 -1 2905
box -2 -3 34 103
use AOI21X1  AOI21X1_131
timestamp 1696145522
transform 1 0 1820 0 -1 2905
box -2 -3 34 103
use AOI21X1  AOI21X1_173
timestamp 1696145522
transform 1 0 1852 0 -1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_174
timestamp 1696145522
transform 1 0 1884 0 -1 2905
box -2 -3 26 103
use INVX1  INVX1_162
timestamp 1696145522
transform 1 0 1908 0 -1 2905
box -2 -3 18 103
use NAND2X1  NAND2X1_306
timestamp 1696145522
transform 1 0 1924 0 -1 2905
box -2 -3 26 103
use NOR2X1  NOR2X1_153
timestamp 1696145522
transform 1 0 1948 0 -1 2905
box -2 -3 26 103
use OAI22X1  OAI22X1_5
timestamp 1696145522
transform -1 0 2012 0 -1 2905
box -2 -3 42 103
use FILL  FILL_28_3_0
timestamp 1696145522
transform 1 0 2012 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_3_1
timestamp 1696145522
transform 1 0 2020 0 -1 2905
box -2 -3 10 103
use AOI22X1  AOI22X1_8
timestamp 1696145522
transform 1 0 2028 0 -1 2905
box -2 -3 42 103
use OAI21X1  OAI21X1_316
timestamp 1696145522
transform -1 0 2100 0 -1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_324
timestamp 1696145522
transform 1 0 2100 0 -1 2905
box -2 -3 26 103
use OR2X2  OR2X2_11
timestamp 1696145522
transform -1 0 2156 0 -1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_546
timestamp 1696145522
transform 1 0 2156 0 -1 2905
box -2 -3 26 103
use NOR2X1  NOR2X1_169
timestamp 1696145522
transform -1 0 2204 0 -1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_327
timestamp 1696145522
transform 1 0 2204 0 -1 2905
box -2 -3 34 103
use INVX2  INVX2_63
timestamp 1696145522
transform 1 0 2236 0 -1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_330
timestamp 1696145522
transform 1 0 2252 0 -1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_154
timestamp 1696145522
transform 1 0 2284 0 -1 2905
box -2 -3 26 103
use NAND3X1  NAND3X1_16
timestamp 1696145522
transform -1 0 2340 0 -1 2905
box -2 -3 34 103
use INVX4  INVX4_19
timestamp 1696145522
transform 1 0 2340 0 -1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_344
timestamp 1696145522
transform -1 0 2388 0 -1 2905
box -2 -3 26 103
use AOI21X1  AOI21X1_89
timestamp 1696145522
transform -1 0 2420 0 -1 2905
box -2 -3 34 103
use AOI21X1  AOI21X1_90
timestamp 1696145522
transform 1 0 2420 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_307
timestamp 1696145522
transform 1 0 2452 0 -1 2905
box -2 -3 34 103
use INVX2  INVX2_64
timestamp 1696145522
transform -1 0 2500 0 -1 2905
box -2 -3 18 103
use AOI21X1  AOI21X1_83
timestamp 1696145522
transform 1 0 2500 0 -1 2905
box -2 -3 34 103
use FILL  FILL_28_4_0
timestamp 1696145522
transform 1 0 2532 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_4_1
timestamp 1696145522
transform 1 0 2540 0 -1 2905
box -2 -3 10 103
use OAI21X1  OAI21X1_285
timestamp 1696145522
transform 1 0 2548 0 -1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_399
timestamp 1696145522
transform -1 0 2604 0 -1 2905
box -2 -3 26 103
use AOI21X1  AOI21X1_96
timestamp 1696145522
transform 1 0 2604 0 -1 2905
box -2 -3 34 103
use OR2X2  OR2X2_9
timestamp 1696145522
transform 1 0 2636 0 -1 2905
box -2 -3 34 103
use NAND3X1  NAND3X1_9
timestamp 1696145522
transform -1 0 2700 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_244
timestamp 1696145522
transform -1 0 2732 0 -1 2905
box -2 -3 34 103
use AND2X2  AND2X2_13
timestamp 1696145522
transform 1 0 2732 0 -1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_135
timestamp 1696145522
transform 1 0 2764 0 -1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_267
timestamp 1696145522
transform 1 0 2788 0 -1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_283
timestamp 1696145522
transform -1 0 2844 0 -1 2905
box -2 -3 34 103
use AND2X2  AND2X2_12
timestamp 1696145522
transform 1 0 2844 0 -1 2905
box -2 -3 34 103
use INVX4  INVX4_17
timestamp 1696145522
transform 1 0 2876 0 -1 2905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_33
timestamp 1696145522
transform 1 0 2900 0 -1 2905
box -2 -3 98 103
use NAND2X1  NAND2X1_138
timestamp 1696145522
transform 1 0 2996 0 -1 2905
box -2 -3 26 103
use INVX1  INVX1_75
timestamp 1696145522
transform -1 0 3036 0 -1 2905
box -2 -3 18 103
use FILL  FILL_28_5_0
timestamp 1696145522
transform 1 0 3036 0 -1 2905
box -2 -3 10 103
use FILL  FILL_28_5_1
timestamp 1696145522
transform 1 0 3044 0 -1 2905
box -2 -3 10 103
use AND2X2  AND2X2_6
timestamp 1696145522
transform 1 0 3052 0 -1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_415
timestamp 1696145522
transform -1 0 3108 0 -1 2905
box -2 -3 26 103
use INVX2  INVX2_51
timestamp 1696145522
transform -1 0 3124 0 -1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_165
timestamp 1696145522
transform 1 0 3124 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_166
timestamp 1696145522
transform -1 0 3188 0 -1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_123
timestamp 1696145522
transform 1 0 3188 0 -1 2905
box -2 -3 26 103
use AOI21X1  AOI21X1_59
timestamp 1696145522
transform 1 0 3212 0 -1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_96
timestamp 1696145522
transform -1 0 3268 0 -1 2905
box -2 -3 26 103
use INVX4  INVX4_1
timestamp 1696145522
transform 1 0 3268 0 -1 2905
box -2 -3 26 103
use AOI21X1  AOI21X1_17
timestamp 1696145522
transform 1 0 3292 0 -1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_35
timestamp 1696145522
transform 1 0 3324 0 -1 2905
box -2 -3 34 103
use AOI21X1  AOI21X1_35
timestamp 1696145522
transform 1 0 3356 0 -1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_91
timestamp 1696145522
transform 1 0 3388 0 -1 2905
box -2 -3 26 103
use AOI21X1  AOI21X1_410
timestamp 1696145522
transform 1 0 3412 0 -1 2905
box -2 -3 34 103
use AOI21X1  AOI21X1_411
timestamp 1696145522
transform -1 0 3476 0 -1 2905
box -2 -3 34 103
use INVX1  INVX1_4
timestamp 1696145522
transform -1 0 3492 0 -1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_943
timestamp 1696145522
transform 1 0 3492 0 -1 2905
box -2 -3 34 103
use AOI21X1  AOI21X1_414
timestamp 1696145522
transform -1 0 3556 0 -1 2905
box -2 -3 34 103
use FILL  FILL_29_1
timestamp 1696145522
transform -1 0 3564 0 -1 2905
box -2 -3 10 103
use AOI21X1  AOI21X1_287
timestamp 1696145522
transform -1 0 36 0 1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_417
timestamp 1696145522
transform 1 0 36 0 1 2905
box -2 -3 26 103
use NOR2X1  NOR2X1_327
timestamp 1696145522
transform 1 0 60 0 1 2905
box -2 -3 26 103
use AOI21X1  AOI21X1_250
timestamp 1696145522
transform 1 0 84 0 1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_339
timestamp 1696145522
transform 1 0 116 0 1 2905
box -2 -3 26 103
use NOR2X1  NOR2X1_328
timestamp 1696145522
transform 1 0 140 0 1 2905
box -2 -3 26 103
use NOR2X1  NOR2X1_329
timestamp 1696145522
transform -1 0 188 0 1 2905
box -2 -3 26 103
use NOR2X1  NOR2X1_348
timestamp 1696145522
transform -1 0 212 0 1 2905
box -2 -3 26 103
use INVX1  INVX1_244
timestamp 1696145522
transform 1 0 212 0 1 2905
box -2 -3 18 103
use AOI22X1  AOI22X1_27
timestamp 1696145522
transform -1 0 268 0 1 2905
box -2 -3 42 103
use OAI21X1  OAI21X1_582
timestamp 1696145522
transform -1 0 300 0 1 2905
box -2 -3 34 103
use INVX1  INVX1_239
timestamp 1696145522
transform -1 0 316 0 1 2905
box -2 -3 18 103
use NOR2X1  NOR2X1_330
timestamp 1696145522
transform -1 0 340 0 1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_572
timestamp 1696145522
transform 1 0 340 0 1 2905
box -2 -3 34 103
use AOI21X1  AOI21X1_224
timestamp 1696145522
transform 1 0 372 0 1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_321
timestamp 1696145522
transform 1 0 404 0 1 2905
box -2 -3 26 103
use NOR2X1  NOR2X1_308
timestamp 1696145522
transform 1 0 428 0 1 2905
box -2 -3 26 103
use NOR2X1  NOR2X1_357
timestamp 1696145522
transform 1 0 452 0 1 2905
box -2 -3 26 103
use INVX1  INVX1_232
timestamp 1696145522
transform 1 0 476 0 1 2905
box -2 -3 18 103
use FILL  FILL_29_0_0
timestamp 1696145522
transform 1 0 492 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_0_1
timestamp 1696145522
transform 1 0 500 0 1 2905
box -2 -3 10 103
use OAI21X1  OAI21X1_564
timestamp 1696145522
transform 1 0 508 0 1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_309
timestamp 1696145522
transform -1 0 564 0 1 2905
box -2 -3 26 103
use NOR2X1  NOR2X1_347
timestamp 1696145522
transform -1 0 588 0 1 2905
box -2 -3 26 103
use INVX2  INVX2_38
timestamp 1696145522
transform 1 0 588 0 1 2905
box -2 -3 18 103
use NOR2X1  NOR2X1_296
timestamp 1696145522
transform 1 0 604 0 1 2905
box -2 -3 26 103
use AND2X2  AND2X2_35
timestamp 1696145522
transform 1 0 628 0 1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_297
timestamp 1696145522
transform -1 0 684 0 1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_660
timestamp 1696145522
transform -1 0 716 0 1 2905
box -2 -3 34 103
use AOI21X1  AOI21X1_288
timestamp 1696145522
transform -1 0 748 0 1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_492
timestamp 1696145522
transform 1 0 748 0 1 2905
box -2 -3 26 103
use INVX1  INVX1_226
timestamp 1696145522
transform 1 0 772 0 1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_662
timestamp 1696145522
transform -1 0 820 0 1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_489
timestamp 1696145522
transform 1 0 820 0 1 2905
box -2 -3 26 103
use AOI22X1  AOI22X1_22
timestamp 1696145522
transform -1 0 884 0 1 2905
box -2 -3 42 103
use INVX1  INVX1_224
timestamp 1696145522
transform 1 0 884 0 1 2905
box -2 -3 18 103
use NOR2X1  NOR2X1_291
timestamp 1696145522
transform 1 0 900 0 1 2905
box -2 -3 26 103
use INVX1  INVX1_229
timestamp 1696145522
transform 1 0 924 0 1 2905
box -2 -3 18 103
use AOI21X1  AOI21X1_216
timestamp 1696145522
transform 1 0 940 0 1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_314
timestamp 1696145522
transform 1 0 972 0 1 2905
box -2 -3 26 103
use FILL  FILL_29_1_0
timestamp 1696145522
transform -1 0 1004 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_1_1
timestamp 1696145522
transform -1 0 1012 0 1 2905
box -2 -3 10 103
use AOI22X1  AOI22X1_23
timestamp 1696145522
transform -1 0 1052 0 1 2905
box -2 -3 42 103
use NOR2X1  NOR2X1_312
timestamp 1696145522
transform 1 0 1052 0 1 2905
box -2 -3 26 103
use NOR2X1  NOR2X1_311
timestamp 1696145522
transform 1 0 1076 0 1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_521
timestamp 1696145522
transform -1 0 1132 0 1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_462
timestamp 1696145522
transform -1 0 1156 0 1 2905
box -2 -3 26 103
use AOI21X1  AOI21X1_192
timestamp 1696145522
transform 1 0 1156 0 1 2905
box -2 -3 34 103
use AOI22X1  AOI22X1_30
timestamp 1696145522
transform 1 0 1188 0 1 2905
box -2 -3 42 103
use NOR2X1  NOR2X1_269
timestamp 1696145522
transform 1 0 1228 0 1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_520
timestamp 1696145522
transform -1 0 1284 0 1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_453
timestamp 1696145522
transform -1 0 1308 0 1 2905
box -2 -3 26 103
use NOR2X1  NOR2X1_281
timestamp 1696145522
transform -1 0 1332 0 1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_659
timestamp 1696145522
transform -1 0 1364 0 1 2905
box -2 -3 34 103
use INVX1  INVX1_203
timestamp 1696145522
transform -1 0 1380 0 1 2905
box -2 -3 18 103
use NAND2X1  NAND2X1_450
timestamp 1696145522
transform -1 0 1404 0 1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_501
timestamp 1696145522
transform -1 0 1436 0 1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_542
timestamp 1696145522
transform -1 0 1460 0 1 2905
box -2 -3 26 103
use NOR2X1  NOR2X1_242
timestamp 1696145522
transform 1 0 1460 0 1 2905
box -2 -3 26 103
use INVX1  INVX1_197
timestamp 1696145522
transform -1 0 1500 0 1 2905
box -2 -3 18 103
use NAND2X1  NAND2X1_443
timestamp 1696145522
transform -1 0 1524 0 1 2905
box -2 -3 26 103
use FILL  FILL_29_2_0
timestamp 1696145522
transform -1 0 1532 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_2_1
timestamp 1696145522
transform -1 0 1540 0 1 2905
box -2 -3 10 103
use OAI21X1  OAI21X1_510
timestamp 1696145522
transform -1 0 1572 0 1 2905
box -2 -3 34 103
use INVX4  INVX4_23
timestamp 1696145522
transform 1 0 1572 0 1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_489
timestamp 1696145522
transform -1 0 1628 0 1 2905
box -2 -3 34 103
use XNOR2X1  XNOR2X1_38
timestamp 1696145522
transform -1 0 1684 0 1 2905
box -2 -3 58 103
use NOR2X1  NOR2X1_241
timestamp 1696145522
transform 1 0 1684 0 1 2905
box -2 -3 26 103
use NOR2X1  NOR2X1_243
timestamp 1696145522
transform 1 0 1708 0 1 2905
box -2 -3 26 103
use OAI22X1  OAI22X1_9
timestamp 1696145522
transform -1 0 1772 0 1 2905
box -2 -3 42 103
use AOI21X1  AOI21X1_189
timestamp 1696145522
transform 1 0 1772 0 1 2905
box -2 -3 34 103
use AOI21X1  AOI21X1_182
timestamp 1696145522
transform -1 0 1836 0 1 2905
box -2 -3 34 103
use AOI21X1  AOI21X1_167
timestamp 1696145522
transform 1 0 1836 0 1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_478
timestamp 1696145522
transform 1 0 1868 0 1 2905
box -2 -3 34 103
use AND2X2  AND2X2_28
timestamp 1696145522
transform -1 0 1932 0 1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_361
timestamp 1696145522
transform -1 0 1964 0 1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_354
timestamp 1696145522
transform 1 0 1964 0 1 2905
box -2 -3 26 103
use AOI21X1  AOI21X1_104
timestamp 1696145522
transform -1 0 2020 0 1 2905
box -2 -3 34 103
use FILL  FILL_29_3_0
timestamp 1696145522
transform -1 0 2028 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_3_1
timestamp 1696145522
transform -1 0 2036 0 1 2905
box -2 -3 10 103
use NAND2X1  NAND2X1_355
timestamp 1696145522
transform -1 0 2060 0 1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_354
timestamp 1696145522
transform -1 0 2092 0 1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_379
timestamp 1696145522
transform 1 0 2092 0 1 2905
box -2 -3 34 103
use AOI21X1  AOI21X1_119
timestamp 1696145522
transform 1 0 2124 0 1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_334
timestamp 1696145522
transform -1 0 2188 0 1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_335
timestamp 1696145522
transform -1 0 2220 0 1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_323
timestamp 1696145522
transform -1 0 2244 0 1 2905
box -2 -3 26 103
use AOI21X1  AOI21X1_111
timestamp 1696145522
transform -1 0 2276 0 1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_181
timestamp 1696145522
transform 1 0 2276 0 1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_363
timestamp 1696145522
transform -1 0 2324 0 1 2905
box -2 -3 26 103
use INVX1  INVX1_142
timestamp 1696145522
transform 1 0 2324 0 1 2905
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_43
timestamp 1696145522
transform 1 0 2340 0 1 2905
box -2 -3 98 103
use NOR2X1  NOR2X1_207
timestamp 1696145522
transform -1 0 2460 0 1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_328
timestamp 1696145522
transform -1 0 2492 0 1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_237
timestamp 1696145522
transform 1 0 2492 0 1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_305
timestamp 1696145522
transform 1 0 2516 0 1 2905
box -2 -3 34 103
use FILL  FILL_29_4_0
timestamp 1696145522
transform -1 0 2556 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_4_1
timestamp 1696145522
transform -1 0 2564 0 1 2905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_48
timestamp 1696145522
transform -1 0 2660 0 1 2905
box -2 -3 98 103
use NOR2X1  NOR2X1_215
timestamp 1696145522
transform 1 0 2660 0 1 2905
box -2 -3 26 103
use NOR2X1  NOR2X1_163
timestamp 1696145522
transform 1 0 2684 0 1 2905
box -2 -3 26 103
use BUFX4  BUFX4_28
timestamp 1696145522
transform -1 0 2740 0 1 2905
box -2 -3 34 103
use CLKBUF1  CLKBUF1_8
timestamp 1696145522
transform -1 0 2812 0 1 2905
box -2 -3 74 103
use INVX2  INVX2_59
timestamp 1696145522
transform 1 0 2812 0 1 2905
box -2 -3 18 103
use OAI21X1  OAI21X1_241
timestamp 1696145522
transform -1 0 2860 0 1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_136
timestamp 1696145522
transform 1 0 2860 0 1 2905
box -2 -3 26 103
use NOR2X1  NOR2X1_144
timestamp 1696145522
transform 1 0 2884 0 1 2905
box -2 -3 26 103
use AOI21X1  AOI21X1_77
timestamp 1696145522
transform 1 0 2908 0 1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_263
timestamp 1696145522
transform 1 0 2940 0 1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_378
timestamp 1696145522
transform 1 0 2972 0 1 2905
box -2 -3 34 103
use NAND2X1  NAND2X1_375
timestamp 1696145522
transform -1 0 3028 0 1 2905
box -2 -3 26 103
use NAND2X1  NAND2X1_139
timestamp 1696145522
transform 1 0 3028 0 1 2905
box -2 -3 26 103
use FILL  FILL_29_5_0
timestamp 1696145522
transform 1 0 3052 0 1 2905
box -2 -3 10 103
use FILL  FILL_29_5_1
timestamp 1696145522
transform 1 0 3060 0 1 2905
box -2 -3 10 103
use NAND2X1  NAND2X1_137
timestamp 1696145522
transform 1 0 3068 0 1 2905
box -2 -3 26 103
use AOI21X1  AOI21X1_39
timestamp 1696145522
transform -1 0 3124 0 1 2905
box -2 -3 34 103
use AOI21X1  AOI21X1_43
timestamp 1696145522
transform -1 0 3156 0 1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_97
timestamp 1696145522
transform 1 0 3156 0 1 2905
box -2 -3 26 103
use OAI21X1  OAI21X1_94
timestamp 1696145522
transform -1 0 3212 0 1 2905
box -2 -3 34 103
use OAI21X1  OAI21X1_93
timestamp 1696145522
transform 1 0 3212 0 1 2905
box -2 -3 34 103
use AOI21X1  AOI21X1_38
timestamp 1696145522
transform 1 0 3244 0 1 2905
box -2 -3 34 103
use BUFX4  BUFX4_29
timestamp 1696145522
transform 1 0 3276 0 1 2905
box -2 -3 34 103
use NOR2X1  NOR2X1_94
timestamp 1696145522
transform 1 0 3308 0 1 2905
box -2 -3 26 103
use NOR2X1  NOR2X1_46
timestamp 1696145522
transform -1 0 3356 0 1 2905
box -2 -3 26 103
use NOR2X1  NOR2X1_47
timestamp 1696145522
transform -1 0 3380 0 1 2905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_29
timestamp 1696145522
transform 1 0 3380 0 1 2905
box -2 -3 98 103
use NOR2X1  NOR2X1_507
timestamp 1696145522
transform -1 0 3500 0 1 2905
box -2 -3 26 103
use NOR2X1  NOR2X1_511
timestamp 1696145522
transform 1 0 3500 0 1 2905
box -2 -3 26 103
use NOR2X1  NOR2X1_404
timestamp 1696145522
transform 1 0 3524 0 1 2905
box -2 -3 26 103
use FILL  FILL_30_1
timestamp 1696145522
transform 1 0 3548 0 1 2905
box -2 -3 10 103
use FILL  FILL_30_2
timestamp 1696145522
transform 1 0 3556 0 1 2905
box -2 -3 10 103
use NOR2X1  NOR2X1_341
timestamp 1696145522
transform -1 0 60 0 1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_589
timestamp 1696145522
transform 1 0 4 0 1 3105
box -2 -3 34 103
use INVX2  INVX2_83
timestamp 1696145522
transform 1 0 28 0 -1 3105
box -2 -3 18 103
use NOR2X1  NOR2X1_340
timestamp 1696145522
transform 1 0 4 0 -1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_506
timestamp 1696145522
transform -1 0 84 0 1 3105
box -2 -3 26 103
use NOR2X1  NOR2X1_332
timestamp 1696145522
transform -1 0 84 0 -1 3105
box -2 -3 26 103
use INVX2  INVX2_86
timestamp 1696145522
transform -1 0 60 0 -1 3105
box -2 -3 18 103
use NAND3X1  NAND3X1_35
timestamp 1696145522
transform -1 0 116 0 1 3105
box -2 -3 34 103
use AND2X2  AND2X2_41
timestamp 1696145522
transform 1 0 108 0 -1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_331
timestamp 1696145522
transform 1 0 84 0 -1 3105
box -2 -3 26 103
use AOI21X1  AOI21X1_245
timestamp 1696145522
transform 1 0 148 0 1 3105
box -2 -3 34 103
use OR2X2  OR2X2_34
timestamp 1696145522
transform -1 0 148 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_590
timestamp 1696145522
transform 1 0 140 0 -1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_240
timestamp 1696145522
transform 1 0 180 0 1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_507
timestamp 1696145522
transform 1 0 172 0 -1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_583
timestamp 1696145522
transform 1 0 244 0 -1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_233
timestamp 1696145522
transform 1 0 212 0 -1 3105
box -2 -3 34 103
use INVX2  INVX2_84
timestamp 1696145522
transform 1 0 196 0 -1 3105
box -2 -3 18 103
use NOR2X1  NOR2X1_326
timestamp 1696145522
transform -1 0 364 0 1 3105
box -2 -3 26 103
use AOI21X1  AOI21X1_231
timestamp 1696145522
transform 1 0 308 0 1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_363
timestamp 1696145522
transform -1 0 388 0 -1 3105
box -2 -3 26 103
use AOI21X1  AOI21X1_238
timestamp 1696145522
transform 1 0 332 0 -1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_335
timestamp 1696145522
transform -1 0 332 0 -1 3105
box -2 -3 26 103
use AOI21X1  AOI21X1_239
timestamp 1696145522
transform 1 0 276 0 -1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_62
timestamp 1696145522
transform -1 0 460 0 1 3105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_59
timestamp 1696145522
transform -1 0 308 0 1 3105
box -2 -3 98 103
use AOI21X1  AOI21X1_258
timestamp 1696145522
transform 1 0 452 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_608
timestamp 1696145522
transform -1 0 452 0 -1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_263
timestamp 1696145522
transform -1 0 420 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_546
timestamp 1696145522
transform 1 0 540 0 1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_283
timestamp 1696145522
transform -1 0 540 0 1 3105
box -2 -3 26 103
use INVX1  INVX1_218
timestamp 1696145522
transform 1 0 500 0 1 3105
box -2 -3 18 103
use FILL  FILL_31_0_1
timestamp 1696145522
transform 1 0 492 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_0_0
timestamp 1696145522
transform 1 0 484 0 1 3105
box -2 -3 10 103
use NOR2X1  NOR2X1_353
timestamp 1696145522
transform 1 0 460 0 1 3105
box -2 -3 26 103
use FILL  FILL_30_0_1
timestamp 1696145522
transform -1 0 500 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_0_0
timestamp 1696145522
transform -1 0 492 0 -1 3105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_61
timestamp 1696145522
transform -1 0 596 0 -1 3105
box -2 -3 98 103
use OAI21X1  OAI21X1_545
timestamp 1696145522
transform 1 0 572 0 1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_284
timestamp 1696145522
transform -1 0 628 0 1 3105
box -2 -3 26 103
use AOI21X1  AOI21X1_257
timestamp 1696145522
transform -1 0 628 0 -1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_545
timestamp 1696145522
transform 1 0 652 0 1 3105
box -2 -3 26 103
use NOR2X1  NOR2X1_293
timestamp 1696145522
transform -1 0 652 0 1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_661
timestamp 1696145522
transform -1 0 684 0 -1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_544
timestamp 1696145522
transform -1 0 652 0 -1 3105
box -2 -3 26 103
use NOR2X1  NOR2X1_285
timestamp 1696145522
transform -1 0 700 0 1 3105
box -2 -3 26 103
use AND2X2  AND2X2_33
timestamp 1696145522
transform 1 0 684 0 -1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_199
timestamp 1696145522
transform -1 0 748 0 1 3105
box -2 -3 34 103
use INVX1  INVX1_223
timestamp 1696145522
transform 1 0 700 0 1 3105
box -2 -3 18 103
use INVX1  INVX1_222
timestamp 1696145522
transform 1 0 716 0 -1 3105
box -2 -3 18 103
use NOR2X1  NOR2X1_276
timestamp 1696145522
transform 1 0 748 0 1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_490
timestamp 1696145522
transform 1 0 756 0 -1 3105
box -2 -3 26 103
use NOR2X1  NOR2X1_310
timestamp 1696145522
transform 1 0 732 0 -1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_533
timestamp 1696145522
transform 1 0 772 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_553
timestamp 1696145522
transform -1 0 812 0 -1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_277
timestamp 1696145522
transform -1 0 860 0 1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_532
timestamp 1696145522
transform 1 0 804 0 1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_201
timestamp 1696145522
transform -1 0 844 0 -1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_476
timestamp 1696145522
transform 1 0 860 0 1 3105
box -2 -3 26 103
use INVX1  INVX1_225
timestamp 1696145522
transform 1 0 868 0 -1 3105
box -2 -3 18 103
use NOR2X1  NOR2X1_292
timestamp 1696145522
transform -1 0 868 0 -1 3105
box -2 -3 26 103
use AOI21X1  AOI21X1_207
timestamp 1696145522
transform 1 0 884 0 1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_202
timestamp 1696145522
transform 1 0 884 0 -1 3105
box -2 -3 34 103
use FILL  FILL_31_1_0
timestamp 1696145522
transform 1 0 996 0 1 3105
box -2 -3 10 103
use NOR2X1  NOR2X1_279
timestamp 1696145522
transform -1 0 996 0 1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_475
timestamp 1696145522
transform -1 0 972 0 1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_543
timestamp 1696145522
transform -1 0 948 0 1 3105
box -2 -3 34 103
use FILL  FILL_30_1_0
timestamp 1696145522
transform -1 0 1004 0 -1 3105
box -2 -3 10 103
use OAI21X1  OAI21X1_563
timestamp 1696145522
transform 1 0 964 0 -1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_307
timestamp 1696145522
transform -1 0 964 0 -1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_486
timestamp 1696145522
transform -1 0 940 0 -1 3105
box -2 -3 26 103
use FILL  FILL_31_1_1
timestamp 1696145522
transform 1 0 1004 0 1 3105
box -2 -3 10 103
use NAND2X1  NAND2X1_488
timestamp 1696145522
transform 1 0 1076 0 -1 3105
box -2 -3 26 103
use INVX2  INVX2_78
timestamp 1696145522
transform -1 0 1076 0 -1 3105
box -2 -3 18 103
use INVX2  INVX2_79
timestamp 1696145522
transform 1 0 1044 0 -1 3105
box -2 -3 18 103
use AND2X2  AND2X2_36
timestamp 1696145522
transform -1 0 1044 0 -1 3105
box -2 -3 34 103
use FILL  FILL_30_1_1
timestamp 1696145522
transform -1 0 1012 0 -1 3105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_63
timestamp 1696145522
transform 1 0 1012 0 1 3105
box -2 -3 98 103
use AOI21X1  AOI21X1_193
timestamp 1696145522
transform 1 0 1124 0 1 3105
box -2 -3 34 103
use INVX1  INVX1_219
timestamp 1696145522
transform -1 0 1124 0 1 3105
box -2 -3 18 103
use AOI21X1  AOI21X1_211
timestamp 1696145522
transform 1 0 1124 0 -1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_487
timestamp 1696145522
transform 1 0 1100 0 -1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_522
timestamp 1696145522
transform 1 0 1156 0 1 3105
box -2 -3 34 103
use OR2X2  OR2X2_33
timestamp 1696145522
transform 1 0 1156 0 -1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_519
timestamp 1696145522
transform -1 0 1220 0 1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_214
timestamp 1696145522
transform 1 0 1188 0 -1 3105
box -2 -3 34 103
use NAND3X1  NAND3X1_31
timestamp 1696145522
transform 1 0 1236 0 1 3105
box -2 -3 34 103
use INVX1  INVX1_216
timestamp 1696145522
transform -1 0 1236 0 1 3105
box -2 -3 18 103
use AOI21X1  AOI21X1_191
timestamp 1696145522
transform -1 0 1252 0 -1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_463
timestamp 1696145522
transform 1 0 1268 0 1 3105
box -2 -3 26 103
use NOR2X1  NOR2X1_278
timestamp 1696145522
transform 1 0 1252 0 -1 3105
box -2 -3 26 103
use XNOR2X1  XNOR2X1_39
timestamp 1696145522
transform -1 0 1348 0 1 3105
box -2 -3 58 103
use NAND2X1  NAND2X1_460
timestamp 1696145522
transform -1 0 1348 0 -1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_518
timestamp 1696145522
transform -1 0 1324 0 -1 3105
box -2 -3 34 103
use INVX2  INVX2_76
timestamp 1696145522
transform -1 0 1292 0 -1 3105
box -2 -3 18 103
use AOI21X1  AOI21X1_197
timestamp 1696145522
transform 1 0 1372 0 1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_257
timestamp 1696145522
transform -1 0 1372 0 1 3105
box -2 -3 26 103
use NOR2X1  NOR2X1_261
timestamp 1696145522
transform -1 0 1396 0 -1 3105
box -2 -3 26 103
use NOR2X1  NOR2X1_258
timestamp 1696145522
transform 1 0 1348 0 -1 3105
box -2 -3 26 103
use AOI21X1  AOI21X1_176
timestamp 1696145522
transform -1 0 1452 0 1 3105
box -2 -3 34 103
use INVX1  INVX1_208
timestamp 1696145522
transform 1 0 1404 0 1 3105
box -2 -3 18 103
use NOR2X1  NOR2X1_263
timestamp 1696145522
transform -1 0 1452 0 -1 3105
box -2 -3 26 103
use AOI21X1  AOI21X1_175
timestamp 1696145522
transform -1 0 1428 0 -1 3105
box -2 -3 34 103
use FILL  FILL_31_2_1
timestamp 1696145522
transform 1 0 1476 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_2_0
timestamp 1696145522
transform 1 0 1468 0 1 3105
box -2 -3 10 103
use INVX1  INVX1_207
timestamp 1696145522
transform -1 0 1468 0 1 3105
box -2 -3 18 103
use NOR2X1  NOR2X1_272
timestamp 1696145522
transform -1 0 1548 0 -1 3105
box -2 -3 26 103
use FILL  FILL_30_2_1
timestamp 1696145522
transform -1 0 1524 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_2_0
timestamp 1696145522
transform -1 0 1516 0 -1 3105
box -2 -3 10 103
use AOI21X1  AOI21X1_223
timestamp 1696145522
transform 1 0 1476 0 -1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_449
timestamp 1696145522
transform -1 0 1476 0 -1 3105
box -2 -3 26 103
use XNOR2X1  XNOR2X1_37
timestamp 1696145522
transform 1 0 1604 0 1 3105
box -2 -3 58 103
use NOR2X1  NOR2X1_303
timestamp 1696145522
transform -1 0 1604 0 1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_509
timestamp 1696145522
transform 1 0 1620 0 -1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_186
timestamp 1696145522
transform 1 0 1588 0 -1 3105
box -2 -3 34 103
use INVX1  INVX1_212
timestamp 1696145522
transform -1 0 1588 0 -1 3105
box -2 -3 18 103
use NOR2X1  NOR2X1_273
timestamp 1696145522
transform -1 0 1572 0 -1 3105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_57
timestamp 1696145522
transform 1 0 1484 0 1 3105
box -2 -3 98 103
use INVX1  INVX1_204
timestamp 1696145522
transform 1 0 1660 0 1 3105
box -2 -3 18 103
use AOI21X1  AOI21X1_184
timestamp 1696145522
transform 1 0 1652 0 -1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_171
timestamp 1696145522
transform -1 0 1708 0 1 3105
box -2 -3 34 103
use BUFX4  BUFX4_30
timestamp 1696145522
transform -1 0 1732 0 -1 3105
box -2 -3 34 103
use INVX2  INVX2_66
timestamp 1696145522
transform -1 0 1700 0 -1 3105
box -2 -3 18 103
use NOR2X1  NOR2X1_259
timestamp 1696145522
transform 1 0 1740 0 1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_488
timestamp 1696145522
transform 1 0 1708 0 1 3105
box -2 -3 34 103
use BUFX4  BUFX4_32
timestamp 1696145522
transform 1 0 1732 0 -1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_246
timestamp 1696145522
transform 1 0 1764 0 1 3105
box -2 -3 26 103
use BUFX4  BUFX4_98
timestamp 1696145522
transform -1 0 1796 0 -1 3105
box -2 -3 34 103
use AND2X2  AND2X2_26
timestamp 1696145522
transform -1 0 1820 0 1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_190
timestamp 1696145522
transform 1 0 1796 0 -1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_275
timestamp 1696145522
transform 1 0 1852 0 1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_473
timestamp 1696145522
transform -1 0 1852 0 1 3105
box -2 -3 34 103
use OAI21X1  OAI21X1_360
timestamp 1696145522
transform 1 0 1892 0 -1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_418
timestamp 1696145522
transform -1 0 1892 0 -1 3105
box -2 -3 26 103
use INVX2  INVX2_70
timestamp 1696145522
transform 1 0 1852 0 -1 3105
box -2 -3 18 103
use NAND2X1  NAND2X1_353
timestamp 1696145522
transform 1 0 1828 0 -1 3105
box -2 -3 26 103
use AOI21X1  AOI21X1_174
timestamp 1696145522
transform 1 0 1972 0 1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_109
timestamp 1696145522
transform 1 0 1980 0 -1 3105
box -2 -3 34 103
use XNOR2X1  XNOR2X1_33
timestamp 1696145522
transform 1 0 1924 0 -1 3105
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_52
timestamp 1696145522
transform 1 0 1876 0 1 3105
box -2 -3 98 103
use FILL  FILL_31_3_1
timestamp 1696145522
transform 1 0 2012 0 1 3105
box -2 -3 10 103
use FILL  FILL_31_3_0
timestamp 1696145522
transform 1 0 2004 0 1 3105
box -2 -3 10 103
use AOI21X1  AOI21X1_99
timestamp 1696145522
transform -1 0 2116 0 -1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_103
timestamp 1696145522
transform -1 0 2084 0 -1 3105
box -2 -3 34 103
use FILL  FILL_30_3_1
timestamp 1696145522
transform -1 0 2052 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_3_0
timestamp 1696145522
transform -1 0 2044 0 -1 3105
box -2 -3 10 103
use NOR2X1  NOR2X1_173
timestamp 1696145522
transform -1 0 2036 0 -1 3105
box -2 -3 26 103
use AOI21X1  AOI21X1_290
timestamp 1696145522
transform -1 0 2204 0 1 3105
box -2 -3 34 103
use BUFX4  BUFX4_102
timestamp 1696145522
transform 1 0 2140 0 1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_255
timestamp 1696145522
transform 1 0 2116 0 1 3105
box -2 -3 26 103
use OR2X2  OR2X2_12
timestamp 1696145522
transform 1 0 2148 0 -1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_124
timestamp 1696145522
transform 1 0 2116 0 -1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_50
timestamp 1696145522
transform 1 0 2020 0 1 3105
box -2 -3 98 103
use NAND2X1  NAND2X1_341
timestamp 1696145522
transform 1 0 2252 0 1 3105
box -2 -3 26 103
use NOR2X1  NOR2X1_214
timestamp 1696145522
transform 1 0 2228 0 1 3105
box -2 -3 26 103
use NOR2X1  NOR2X1_419
timestamp 1696145522
transform 1 0 2204 0 1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_357
timestamp 1696145522
transform -1 0 2268 0 -1 3105
box -2 -3 34 103
use INVX1  INVX1_143
timestamp 1696145522
transform -1 0 2236 0 -1 3105
box -2 -3 18 103
use AOI22X1  AOI22X1_9
timestamp 1696145522
transform -1 0 2220 0 -1 3105
box -2 -3 42 103
use OAI21X1  OAI21X1_346
timestamp 1696145522
transform 1 0 2316 0 1 3105
box -2 -3 34 103
use NAND2X1  NAND2X1_342
timestamp 1696145522
transform -1 0 2316 0 1 3105
box -2 -3 26 103
use INVX2  INVX2_67
timestamp 1696145522
transform 1 0 2276 0 1 3105
box -2 -3 18 103
use NAND2X1  NAND2X1_343
timestamp 1696145522
transform 1 0 2268 0 -1 3105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_42
timestamp 1696145522
transform 1 0 2348 0 1 3105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_44
timestamp 1696145522
transform -1 0 2388 0 -1 3105
box -2 -3 98 103
use INVX2  INVX2_68
timestamp 1696145522
transform 1 0 2388 0 -1 3105
box -2 -3 18 103
use NAND2X1  NAND2X1_345
timestamp 1696145522
transform -1 0 2452 0 -1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_356
timestamp 1696145522
transform 1 0 2404 0 -1 3105
box -2 -3 26 103
use NOR2X1  NOR2X1_187
timestamp 1696145522
transform -1 0 2468 0 1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_329
timestamp 1696145522
transform 1 0 2452 0 -1 3105
box -2 -3 34 103
use INVX1  INVX1_148
timestamp 1696145522
transform 1 0 2492 0 1 3105
box -2 -3 18 103
use NOR2X1  NOR2X1_383
timestamp 1696145522
transform 1 0 2468 0 1 3105
box -2 -3 26 103
use AOI21X1  AOI21X1_97
timestamp 1696145522
transform 1 0 2484 0 -1 3105
box -2 -3 34 103
use FILL  FILL_31_4_0
timestamp 1696145522
transform 1 0 2532 0 1 3105
box -2 -3 10 103
use NOR2X1  NOR2X1_236
timestamp 1696145522
transform 1 0 2508 0 1 3105
box -2 -3 26 103
use AOI21X1  AOI21X1_158
timestamp 1696145522
transform 1 0 2516 0 -1 3105
box -2 -3 34 103
use FILL  FILL_31_4_1
timestamp 1696145522
transform 1 0 2540 0 1 3105
box -2 -3 10 103
use OAI21X1  OAI21X1_344
timestamp 1696145522
transform 1 0 2564 0 -1 3105
box -2 -3 34 103
use FILL  FILL_30_4_1
timestamp 1696145522
transform 1 0 2556 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_4_0
timestamp 1696145522
transform 1 0 2548 0 -1 3105
box -2 -3 10 103
use NAND2X1  NAND2X1_531
timestamp 1696145522
transform -1 0 2732 0 1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_347
timestamp 1696145522
transform 1 0 2676 0 1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_102
timestamp 1696145522
transform 1 0 2644 0 1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_47
timestamp 1696145522
transform 1 0 2548 0 1 3105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_38
timestamp 1696145522
transform 1 0 2692 0 -1 3105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_45
timestamp 1696145522
transform 1 0 2596 0 -1 3105
box -2 -3 98 103
use BUFX4  BUFX4_101
timestamp 1696145522
transform -1 0 2820 0 -1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_76
timestamp 1696145522
transform 1 0 2820 0 -1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_143
timestamp 1696145522
transform 1 0 2852 0 -1 3105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_34
timestamp 1696145522
transform 1 0 2876 0 -1 3105
box -2 -3 98 103
use NOR2X1  NOR2X1_382
timestamp 1696145522
transform -1 0 2756 0 1 3105
box -2 -3 26 103
use BUFX2  BUFX2_47
timestamp 1696145522
transform 1 0 2756 0 1 3105
box -2 -3 26 103
use AOI21X1  AOI21X1_110
timestamp 1696145522
transform 1 0 2780 0 1 3105
box -2 -3 34 103
use NOR2X1  NOR2X1_172
timestamp 1696145522
transform 1 0 2812 0 1 3105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_35
timestamp 1696145522
transform 1 0 2836 0 1 3105
box -2 -3 98 103
use NOR2X1  NOR2X1_379
timestamp 1696145522
transform 1 0 2956 0 1 3105
box -2 -3 26 103
use BUFX2  BUFX2_35
timestamp 1696145522
transform -1 0 2956 0 1 3105
box -2 -3 26 103
use NOR2X1  NOR2X1_133
timestamp 1696145522
transform -1 0 2996 0 -1 3105
box -2 -3 26 103
use FILL  FILL_31_5_0
timestamp 1696145522
transform 1 0 3076 0 1 3105
box -2 -3 10 103
use INVX1  INVX1_125
timestamp 1696145522
transform -1 0 3092 0 -1 3105
box -2 -3 18 103
use FILL  FILL_30_5_1
timestamp 1696145522
transform -1 0 3076 0 -1 3105
box -2 -3 10 103
use FILL  FILL_30_5_0
timestamp 1696145522
transform -1 0 3068 0 -1 3105
box -2 -3 10 103
use OAI21X1  OAI21X1_306
timestamp 1696145522
transform 1 0 3028 0 -1 3105
box -2 -3 34 103
use AOI21X1  AOI21X1_81
timestamp 1696145522
transform 1 0 2996 0 -1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_41
timestamp 1696145522
transform 1 0 2980 0 1 3105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_37
timestamp 1696145522
transform 1 0 3092 0 -1 3105
box -2 -3 98 103
use AOI21X1  AOI21X1_44
timestamp 1696145522
transform 1 0 3188 0 -1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_32
timestamp 1696145522
transform 1 0 3220 0 -1 3105
box -2 -3 98 103
use FILL  FILL_31_5_1
timestamp 1696145522
transform 1 0 3084 0 1 3105
box -2 -3 10 103
use NOR2X1  NOR2X1_152
timestamp 1696145522
transform 1 0 3092 0 1 3105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_36
timestamp 1696145522
transform 1 0 3116 0 1 3105
box -2 -3 98 103
use NOR2X1  NOR2X1_377
timestamp 1696145522
transform -1 0 3236 0 1 3105
box -2 -3 26 103
use NOR2X1  NOR2X1_376
timestamp 1696145522
transform 1 0 3236 0 1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_529
timestamp 1696145522
transform 1 0 3260 0 1 3105
box -2 -3 26 103
use NOR2X1  NOR2X1_93
timestamp 1696145522
transform -1 0 3356 0 1 3105
box -2 -3 26 103
use NAND2X1  NAND2X1_530
timestamp 1696145522
transform -1 0 3332 0 1 3105
box -2 -3 26 103
use NOR2X1  NOR2X1_380
timestamp 1696145522
transform 1 0 3284 0 1 3105
box -2 -3 26 103
use OAI21X1  OAI21X1_24
timestamp 1696145522
transform 1 0 3332 0 -1 3105
box -2 -3 34 103
use INVX1  INVX1_26
timestamp 1696145522
transform 1 0 3316 0 -1 3105
box -2 -3 18 103
use NOR2X1  NOR2X1_92
timestamp 1696145522
transform -1 0 3404 0 1 3105
box -2 -3 26 103
use NOR2X1  NOR2X1_378
timestamp 1696145522
transform -1 0 3380 0 1 3105
box -2 -3 26 103
use AOI21X1  AOI21X1_37
timestamp 1696145522
transform 1 0 3364 0 -1 3105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_31
timestamp 1696145522
transform -1 0 3500 0 1 3105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_30
timestamp 1696145522
transform 1 0 3396 0 -1 3105
box -2 -3 98 103
use BUFX2  BUFX2_32
timestamp 1696145522
transform 1 0 3492 0 -1 3105
box -2 -3 26 103
use INVX1  INVX1_273
timestamp 1696145522
transform -1 0 3532 0 -1 3105
box -2 -3 18 103
use BUFX2  BUFX2_31
timestamp 1696145522
transform 1 0 3532 0 -1 3105
box -2 -3 26 103
use FILL  FILL_31_1
timestamp 1696145522
transform -1 0 3564 0 -1 3105
box -2 -3 10 103
use BUFX4  BUFX4_103
timestamp 1696145522
transform -1 0 3532 0 1 3105
box -2 -3 34 103
use BUFX2  BUFX2_23
timestamp 1696145522
transform 1 0 3532 0 1 3105
box -2 -3 26 103
use FILL  FILL_32_1
timestamp 1696145522
transform 1 0 3556 0 1 3105
box -2 -3 10 103
use BUFX2  BUFX2_62
timestamp 1696145522
transform -1 0 28 0 -1 3305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_60
timestamp 1696145522
transform -1 0 124 0 -1 3305
box -2 -3 98 103
use AOI21X1  AOI21X1_246
timestamp 1696145522
transform 1 0 124 0 -1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_336
timestamp 1696145522
transform -1 0 180 0 -1 3305
box -2 -3 26 103
use BUFX2  BUFX2_61
timestamp 1696145522
transform -1 0 204 0 -1 3305
box -2 -3 26 103
use NOR2X1  NOR2X1_392
timestamp 1696145522
transform -1 0 228 0 -1 3305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_58
timestamp 1696145522
transform 1 0 228 0 -1 3305
box -2 -3 98 103
use BUFX2  BUFX2_64
timestamp 1696145522
transform -1 0 348 0 -1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_534
timestamp 1696145522
transform -1 0 372 0 -1 3305
box -2 -3 26 103
use NOR2X1  NOR2X1_391
timestamp 1696145522
transform -1 0 396 0 -1 3305
box -2 -3 26 103
use BUFX2  BUFX2_63
timestamp 1696145522
transform 1 0 396 0 -1 3305
box -2 -3 26 103
use NOR2X1  NOR2X1_393
timestamp 1696145522
transform -1 0 444 0 -1 3305
box -2 -3 26 103
use OR2X2  OR2X2_37
timestamp 1696145522
transform -1 0 476 0 -1 3305
box -2 -3 34 103
use BUFX2  BUFX2_60
timestamp 1696145522
transform 1 0 476 0 -1 3305
box -2 -3 26 103
use FILL  FILL_32_0_0
timestamp 1696145522
transform 1 0 500 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_0_1
timestamp 1696145522
transform 1 0 508 0 -1 3305
box -2 -3 10 103
use BUFX2  BUFX2_57
timestamp 1696145522
transform 1 0 516 0 -1 3305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_55
timestamp 1696145522
transform -1 0 636 0 -1 3305
box -2 -3 98 103
use NOR2X1  NOR2X1_295
timestamp 1696145522
transform -1 0 660 0 -1 3305
box -2 -3 26 103
use AOI21X1  AOI21X1_208
timestamp 1696145522
transform -1 0 692 0 -1 3305
box -2 -3 34 103
use AND2X2  AND2X2_32
timestamp 1696145522
transform 1 0 692 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_544
timestamp 1696145522
transform -1 0 756 0 -1 3305
box -2 -3 34 103
use AOI21X1  AOI21X1_200
timestamp 1696145522
transform 1 0 756 0 -1 3305
box -2 -3 34 103
use CLKBUF1  CLKBUF1_5
timestamp 1696145522
transform -1 0 860 0 -1 3305
box -2 -3 74 103
use AOI21X1  AOI21X1_209
timestamp 1696145522
transform 1 0 860 0 -1 3305
box -2 -3 34 103
use AOI21X1  AOI21X1_210
timestamp 1696145522
transform -1 0 924 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_552
timestamp 1696145522
transform -1 0 956 0 -1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_280
timestamp 1696145522
transform 1 0 956 0 -1 3305
box -2 -3 26 103
use NOR2X1  NOR2X1_286
timestamp 1696145522
transform -1 0 1004 0 -1 3305
box -2 -3 26 103
use FILL  FILL_32_1_0
timestamp 1696145522
transform -1 0 1012 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_1_1
timestamp 1696145522
transform -1 0 1020 0 -1 3305
box -2 -3 10 103
use AOI21X1  AOI21X1_195
timestamp 1696145522
transform -1 0 1052 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_531
timestamp 1696145522
transform -1 0 1084 0 -1 3305
box -2 -3 34 103
use AOI21X1  AOI21X1_215
timestamp 1696145522
transform 1 0 1084 0 -1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_302
timestamp 1696145522
transform 1 0 1116 0 -1 3305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_56
timestamp 1696145522
transform -1 0 1236 0 -1 3305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_54
timestamp 1696145522
transform 1 0 1236 0 -1 3305
box -2 -3 98 103
use AOI21X1  AOI21X1_198
timestamp 1696145522
transform 1 0 1332 0 -1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_289
timestamp 1696145522
transform -1 0 1388 0 -1 3305
box -2 -3 26 103
use CLKBUF1  CLKBUF1_4
timestamp 1696145522
transform -1 0 1460 0 -1 3305
box -2 -3 74 103
use AOI21X1  AOI21X1_177
timestamp 1696145522
transform -1 0 1492 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_498
timestamp 1696145522
transform -1 0 1524 0 -1 3305
box -2 -3 34 103
use FILL  FILL_32_2_0
timestamp 1696145522
transform 1 0 1524 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_2_1
timestamp 1696145522
transform 1 0 1532 0 -1 3305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_51
timestamp 1696145522
transform 1 0 1540 0 -1 3305
box -2 -3 98 103
use AOI21X1  AOI21X1_185
timestamp 1696145522
transform 1 0 1636 0 -1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_260
timestamp 1696145522
transform -1 0 1692 0 -1 3305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_49
timestamp 1696145522
transform 1 0 1692 0 -1 3305
box -2 -3 98 103
use NOR2X1  NOR2X1_240
timestamp 1696145522
transform -1 0 1812 0 -1 3305
box -2 -3 26 103
use AOI21X1  AOI21X1_170
timestamp 1696145522
transform -1 0 1844 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_529
timestamp 1696145522
transform 1 0 1844 0 -1 3305
box -2 -3 34 103
use OAI21X1  OAI21X1_530
timestamp 1696145522
transform -1 0 1908 0 -1 3305
box -2 -3 34 103
use INVX1  INVX1_215
timestamp 1696145522
transform -1 0 1924 0 -1 3305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_53
timestamp 1696145522
transform 1 0 1924 0 -1 3305
box -2 -3 98 103
use FILL  FILL_32_3_0
timestamp 1696145522
transform 1 0 2020 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_3_1
timestamp 1696145522
transform 1 0 2028 0 -1 3305
box -2 -3 10 103
use BUFX2  BUFX2_56
timestamp 1696145522
transform 1 0 2036 0 -1 3305
box -2 -3 26 103
use NOR2X1  NOR2X1_385
timestamp 1696145522
transform -1 0 2084 0 -1 3305
box -2 -3 26 103
use BUFX2  BUFX2_55
timestamp 1696145522
transform 1 0 2084 0 -1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_532
timestamp 1696145522
transform 1 0 2108 0 -1 3305
box -2 -3 26 103
use NOR2X1  NOR2X1_386
timestamp 1696145522
transform -1 0 2156 0 -1 3305
box -2 -3 26 103
use BUFX2  BUFX2_54
timestamp 1696145522
transform 1 0 2156 0 -1 3305
box -2 -3 26 103
use NOR2X1  NOR2X1_390
timestamp 1696145522
transform 1 0 2180 0 -1 3305
box -2 -3 26 103
use NAND3X1  NAND3X1_43
timestamp 1696145522
transform 1 0 2204 0 -1 3305
box -2 -3 34 103
use NOR2X1  NOR2X1_389
timestamp 1696145522
transform 1 0 2236 0 -1 3305
box -2 -3 26 103
use BUFX2  BUFX2_53
timestamp 1696145522
transform 1 0 2260 0 -1 3305
box -2 -3 26 103
use BUFX2  BUFX2_59
timestamp 1696145522
transform 1 0 2284 0 -1 3305
box -2 -3 26 103
use BUFX2  BUFX2_58
timestamp 1696145522
transform 1 0 2308 0 -1 3305
box -2 -3 26 103
use BUFX2  BUFX2_52
timestamp 1696145522
transform 1 0 2332 0 -1 3305
box -2 -3 26 103
use NOR2X1  NOR2X1_387
timestamp 1696145522
transform -1 0 2380 0 -1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_533
timestamp 1696145522
transform 1 0 2380 0 -1 3305
box -2 -3 26 103
use BUFX2  BUFX2_45
timestamp 1696145522
transform -1 0 2428 0 -1 3305
box -2 -3 26 103
use BUFX2  BUFX2_65
timestamp 1696145522
transform -1 0 2452 0 -1 3305
box -2 -3 26 103
use BUFX2  BUFX2_51
timestamp 1696145522
transform 1 0 2452 0 -1 3305
box -2 -3 26 103
use BUFX2  BUFX2_46
timestamp 1696145522
transform 1 0 2476 0 -1 3305
box -2 -3 26 103
use NOR2X1  NOR2X1_388
timestamp 1696145522
transform -1 0 2524 0 -1 3305
box -2 -3 26 103
use BUFX2  BUFX2_66
timestamp 1696145522
transform 1 0 2524 0 -1 3305
box -2 -3 26 103
use FILL  FILL_32_4_0
timestamp 1696145522
transform 1 0 2548 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_4_1
timestamp 1696145522
transform 1 0 2556 0 -1 3305
box -2 -3 10 103
use BUFX2  BUFX2_50
timestamp 1696145522
transform 1 0 2564 0 -1 3305
box -2 -3 26 103
use BUFX2  BUFX2_49
timestamp 1696145522
transform 1 0 2588 0 -1 3305
box -2 -3 26 103
use BUFX2  BUFX2_44
timestamp 1696145522
transform 1 0 2612 0 -1 3305
box -2 -3 26 103
use OR2X2  OR2X2_36
timestamp 1696145522
transform -1 0 2668 0 -1 3305
box -2 -3 34 103
use BUFX2  BUFX2_48
timestamp 1696145522
transform 1 0 2668 0 -1 3305
box -2 -3 26 103
use NOR2X1  NOR2X1_384
timestamp 1696145522
transform 1 0 2692 0 -1 3305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_40
timestamp 1696145522
transform -1 0 2812 0 -1 3305
box -2 -3 98 103
use INVX1  INVX1_141
timestamp 1696145522
transform 1 0 2812 0 -1 3305
box -2 -3 18 103
use OAI21X1  OAI21X1_345
timestamp 1696145522
transform -1 0 2860 0 -1 3305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_39
timestamp 1696145522
transform 1 0 2860 0 -1 3305
box -2 -3 98 103
use BUFX2  BUFX2_36
timestamp 1696145522
transform 1 0 2956 0 -1 3305
box -2 -3 26 103
use BUFX2  BUFX2_41
timestamp 1696145522
transform 1 0 2980 0 -1 3305
box -2 -3 26 103
use BUFX2  BUFX2_43
timestamp 1696145522
transform 1 0 3004 0 -1 3305
box -2 -3 26 103
use BUFX2  BUFX2_42
timestamp 1696145522
transform 1 0 3028 0 -1 3305
box -2 -3 26 103
use FILL  FILL_32_5_0
timestamp 1696145522
transform 1 0 3052 0 -1 3305
box -2 -3 10 103
use FILL  FILL_32_5_1
timestamp 1696145522
transform 1 0 3060 0 -1 3305
box -2 -3 10 103
use NOR2X1  NOR2X1_381
timestamp 1696145522
transform 1 0 3068 0 -1 3305
box -2 -3 26 103
use NOR2X1  NOR2X1_394
timestamp 1696145522
transform -1 0 3116 0 -1 3305
box -2 -3 26 103
use NAND3X1  NAND3X1_42
timestamp 1696145522
transform 1 0 3116 0 -1 3305
box -2 -3 34 103
use BUFX2  BUFX2_40
timestamp 1696145522
transform -1 0 3172 0 -1 3305
box -2 -3 26 103
use BUFX2  BUFX2_39
timestamp 1696145522
transform 1 0 3172 0 -1 3305
box -2 -3 26 103
use BUFX2  BUFX2_38
timestamp 1696145522
transform 1 0 3196 0 -1 3305
box -2 -3 26 103
use BUFX2  BUFX2_37
timestamp 1696145522
transform 1 0 3220 0 -1 3305
box -2 -3 26 103
use CLKBUF1  CLKBUF1_3
timestamp 1696145522
transform -1 0 3316 0 -1 3305
box -2 -3 74 103
use BUFX2  BUFX2_34
timestamp 1696145522
transform -1 0 3340 0 -1 3305
box -2 -3 26 103
use BUFX2  BUFX2_33
timestamp 1696145522
transform -1 0 3364 0 -1 3305
box -2 -3 26 103
use NOR2X1  NOR2X1_48
timestamp 1696145522
transform -1 0 3388 0 -1 3305
box -2 -3 26 103
use OAI21X1  OAI21X1_901
timestamp 1696145522
transform 1 0 3388 0 -1 3305
box -2 -3 34 103
use NAND2X1  NAND2X1_81
timestamp 1696145522
transform -1 0 3444 0 -1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_641
timestamp 1696145522
transform -1 0 3468 0 -1 3305
box -2 -3 26 103
use NAND2X1  NAND2X1_642
timestamp 1696145522
transform -1 0 3492 0 -1 3305
box -2 -3 26 103
use NOR2X1  NOR2X1_407
timestamp 1696145522
transform -1 0 3516 0 -1 3305
box -2 -3 26 103
use AND2X2  AND2X2_45
timestamp 1696145522
transform 1 0 3516 0 -1 3305
box -2 -3 34 103
use FILL  FILL_33_1
timestamp 1696145522
transform -1 0 3556 0 -1 3305
box -2 -3 10 103
use FILL  FILL_33_2
timestamp 1696145522
transform -1 0 3564 0 -1 3305
box -2 -3 10 103
<< labels >>
flabel metal6 s 480 -30 496 -22 7 FreeSans 24 270 0 0 vdd
port 0 nsew
flabel metal6 s 992 -30 1008 -22 7 FreeSans 24 270 0 0 gnd
port 1 nsew
flabel metal2 s 854 3328 858 3332 3 FreeSans 24 90 0 0 clk
port 2 nsew
flabel metal3 s 3590 1728 3594 1732 3 FreeSans 24 0 0 0 reset
port 3 nsew
flabel metal2 s 1214 -22 1218 -18 7 FreeSans 24 270 0 0 operand_A[0]
port 4 nsew
flabel metal2 s 902 -22 906 -18 7 FreeSans 24 270 0 0 operand_A[1]
port 5 nsew
flabel metal2 s 886 -22 890 -18 7 FreeSans 24 270 0 0 operand_A[2]
port 6 nsew
flabel metal2 s 1334 -22 1338 -18 7 FreeSans 24 270 0 0 operand_A[3]
port 7 nsew
flabel metal2 s 1270 -22 1274 -18 7 FreeSans 24 270 0 0 operand_A[4]
port 8 nsew
flabel metal2 s 838 -22 842 -18 7 FreeSans 24 270 0 0 operand_A[5]
port 9 nsew
flabel metal2 s 646 -22 650 -18 7 FreeSans 24 270 0 0 operand_A[6]
port 10 nsew
flabel metal2 s 694 -22 698 -18 7 FreeSans 24 270 0 0 operand_A[7]
port 11 nsew
flabel metal2 s 1070 -22 1074 -18 7 FreeSans 24 270 0 0 operand_A[8]
port 12 nsew
flabel metal2 s 2582 -22 2586 -18 7 FreeSans 24 270 0 0 operand_A[9]
port 13 nsew
flabel metal2 s 518 -22 522 -18 7 FreeSans 24 270 0 0 operand_A[10]
port 14 nsew
flabel metal2 s 622 -22 626 -18 7 FreeSans 24 270 0 0 operand_A[11]
port 15 nsew
flabel metal2 s 982 -22 986 -18 7 FreeSans 24 270 0 0 operand_A[12]
port 16 nsew
flabel metal2 s 782 -22 786 -18 7 FreeSans 24 270 0 0 operand_A[13]
port 17 nsew
flabel metal2 s 806 -22 810 -18 7 FreeSans 24 270 0 0 operand_A[14]
port 18 nsew
flabel metal2 s 2886 -22 2890 -18 7 FreeSans 24 270 0 0 operand_A[15]
port 19 nsew
flabel metal2 s 1046 -22 1050 -18 7 FreeSans 24 270 0 0 operand_A[16]
port 20 nsew
flabel metal2 s 606 -22 610 -18 7 FreeSans 24 270 0 0 operand_A[17]
port 21 nsew
flabel metal3 s 3590 1078 3594 1082 3 FreeSans 24 0 0 0 operand_A[18]
port 22 nsew
flabel metal3 s 3590 888 3594 892 3 FreeSans 24 0 0 0 operand_A[19]
port 23 nsew
flabel metal3 s -26 958 -22 962 7 FreeSans 24 0 0 0 operand_A[20]
port 24 nsew
flabel metal3 s 3590 1348 3594 1352 3 FreeSans 24 0 0 0 operand_A[21]
port 25 nsew
flabel metal3 s 3590 1788 3594 1792 3 FreeSans 24 0 0 0 operand_A[22]
port 26 nsew
flabel metal3 s 3590 1868 3594 1872 3 FreeSans 24 0 0 0 operand_A[23]
port 27 nsew
flabel metal3 s 3590 2148 3594 2152 3 FreeSans 24 0 0 0 operand_A[24]
port 28 nsew
flabel metal3 s 3590 2168 3594 2172 3 FreeSans 24 0 0 0 operand_A[25]
port 29 nsew
flabel metal3 s 3590 2198 3594 2202 3 FreeSans 24 0 0 0 operand_A[26]
port 30 nsew
flabel metal3 s 3590 2258 3594 2262 3 FreeSans 24 0 0 0 operand_A[27]
port 31 nsew
flabel metal3 s 3590 2538 3594 2542 3 FreeSans 24 0 0 0 operand_A[28]
port 32 nsew
flabel metal3 s 3590 2688 3594 2692 3 FreeSans 24 0 0 0 operand_A[29]
port 33 nsew
flabel metal3 s 3590 2728 3594 2732 3 FreeSans 24 0 0 0 operand_A[30]
port 34 nsew
flabel metal2 s 3086 3328 3090 3332 3 FreeSans 24 90 0 0 operand_A[31]
port 35 nsew
flabel metal2 s 2630 3328 2634 3332 3 FreeSans 24 90 0 0 operand_A[32]
port 36 nsew
flabel metal2 s 2526 3328 2530 3332 3 FreeSans 24 90 0 0 operand_A[33]
port 37 nsew
flabel metal2 s 2798 3328 2802 3332 3 FreeSans 24 90 0 0 operand_A[34]
port 38 nsew
flabel metal2 s 2942 3328 2946 3332 3 FreeSans 24 90 0 0 operand_A[35]
port 39 nsew
flabel metal2 s 1950 3328 1954 3332 3 FreeSans 24 90 0 0 operand_A[36]
port 40 nsew
flabel metal2 s 2246 3328 2250 3332 3 FreeSans 24 90 0 0 operand_A[37]
port 41 nsew
flabel metal2 s 2262 3328 2266 3332 3 FreeSans 24 90 0 0 operand_A[38]
port 42 nsew
flabel metal2 s 1886 3328 1890 3332 3 FreeSans 24 90 0 0 operand_A[39]
port 43 nsew
flabel metal2 s 1742 3328 1746 3332 3 FreeSans 24 90 0 0 operand_A[40]
port 44 nsew
flabel metal2 s 1598 3328 1602 3332 3 FreeSans 24 90 0 0 operand_A[41]
port 45 nsew
flabel metal2 s 1054 3328 1058 3332 3 FreeSans 24 90 0 0 operand_A[42]
port 46 nsew
flabel metal3 s -26 2348 -22 2352 7 FreeSans 24 0 0 0 operand_A[43]
port 47 nsew
flabel metal3 s -26 2268 -22 2272 7 FreeSans 24 0 0 0 operand_A[44]
port 48 nsew
flabel metal3 s -26 2248 -22 2252 7 FreeSans 24 0 0 0 operand_A[45]
port 49 nsew
flabel metal2 s 1022 3328 1026 3332 3 FreeSans 24 90 0 0 operand_A[46]
port 50 nsew
flabel metal3 s -26 2368 -22 2372 7 FreeSans 24 0 0 0 operand_A[47]
port 51 nsew
flabel metal2 s 1534 3328 1538 3332 3 FreeSans 24 90 0 0 operand_A[48]
port 52 nsew
flabel metal2 s 1350 3328 1354 3332 3 FreeSans 24 90 0 0 operand_A[49]
port 53 nsew
flabel metal2 s 1390 3328 1394 3332 3 FreeSans 24 90 0 0 operand_A[50]
port 54 nsew
flabel metal2 s 1230 3328 1234 3332 3 FreeSans 24 90 0 0 operand_A[51]
port 55 nsew
flabel metal2 s 710 3328 714 3332 3 FreeSans 24 90 0 0 operand_A[52]
port 56 nsew
flabel metal2 s 606 3328 610 3332 3 FreeSans 24 90 0 0 operand_A[53]
port 57 nsew
flabel metal2 s 694 3328 698 3332 3 FreeSans 24 90 0 0 operand_A[54]
port 58 nsew
flabel metal2 s 630 3328 634 3332 3 FreeSans 24 90 0 0 operand_A[55]
port 59 nsew
flabel metal3 s -26 2398 -22 2402 7 FreeSans 24 0 0 0 operand_A[56]
port 60 nsew
flabel metal3 s -26 2628 -22 2632 7 FreeSans 24 0 0 0 operand_A[57]
port 61 nsew
flabel metal3 s -26 2608 -22 2612 7 FreeSans 24 0 0 0 operand_A[58]
port 62 nsew
flabel metal3 s -26 2848 -22 2852 7 FreeSans 24 0 0 0 operand_A[59]
port 63 nsew
flabel metal3 s -26 2158 -22 2162 7 FreeSans 24 0 0 0 operand_A[60]
port 64 nsew
flabel metal3 s -26 2448 -22 2452 7 FreeSans 24 0 0 0 operand_A[61]
port 65 nsew
flabel metal3 s -26 2178 -22 2182 7 FreeSans 24 0 0 0 operand_A[62]
port 66 nsew
flabel metal3 s -26 2588 -22 2592 7 FreeSans 24 0 0 0 operand_A[63]
port 67 nsew
flabel metal3 s -26 248 -22 252 7 FreeSans 24 0 0 0 operand_B[0]
port 68 nsew
flabel metal2 s 142 -22 146 -18 7 FreeSans 24 270 0 0 operand_B[1]
port 69 nsew
flabel metal3 s -26 348 -22 352 7 FreeSans 24 0 0 0 operand_B[2]
port 70 nsew
flabel metal2 s 286 -22 290 -18 7 FreeSans 24 270 0 0 operand_B[3]
port 71 nsew
flabel metal2 s 1486 -22 1490 -18 7 FreeSans 24 270 0 0 operand_B[4]
port 72 nsew
flabel metal2 s 1542 -22 1546 -18 7 FreeSans 24 270 0 0 operand_B[5]
port 73 nsew
flabel metal2 s 1782 -22 1786 -18 7 FreeSans 24 270 0 0 operand_B[6]
port 74 nsew
flabel metal2 s 1598 -22 1602 -18 7 FreeSans 24 270 0 0 operand_B[7]
port 75 nsew
flabel metal2 s 2206 -22 2210 -18 7 FreeSans 24 270 0 0 operand_B[8]
port 76 nsew
flabel metal2 s 2478 -22 2482 -18 7 FreeSans 24 270 0 0 operand_B[9]
port 77 nsew
flabel metal2 s 3006 -22 3010 -18 7 FreeSans 24 270 0 0 operand_B[10]
port 78 nsew
flabel metal2 s 3150 -22 3154 -18 7 FreeSans 24 270 0 0 operand_B[11]
port 79 nsew
flabel metal2 s 2678 -22 2682 -18 7 FreeSans 24 270 0 0 operand_B[12]
port 80 nsew
flabel metal2 s 2278 -22 2282 -18 7 FreeSans 24 270 0 0 operand_B[13]
port 81 nsew
flabel metal2 s 3350 -22 3354 -18 7 FreeSans 24 270 0 0 operand_B[14]
port 82 nsew
flabel metal2 s 2910 -22 2914 -18 7 FreeSans 24 270 0 0 operand_B[15]
port 83 nsew
flabel metal2 s 2862 -22 2866 -18 7 FreeSans 24 270 0 0 operand_B[16]
port 84 nsew
flabel metal2 s 2702 -22 2706 -18 7 FreeSans 24 270 0 0 operand_B[17]
port 85 nsew
flabel metal3 s 3590 978 3594 982 3 FreeSans 24 0 0 0 operand_B[18]
port 86 nsew
flabel metal3 s 3590 908 3594 912 3 FreeSans 24 0 0 0 operand_B[19]
port 87 nsew
flabel metal3 s 3590 1248 3594 1252 3 FreeSans 24 0 0 0 operand_B[20]
port 88 nsew
flabel metal3 s 3590 1448 3594 1452 3 FreeSans 24 0 0 0 operand_B[21]
port 89 nsew
flabel metal3 s 3590 1768 3594 1772 3 FreeSans 24 0 0 0 operand_B[22]
port 90 nsew
flabel metal3 s 3590 1678 3594 1682 3 FreeSans 24 0 0 0 operand_B[23]
port 91 nsew
flabel metal3 s 3590 2098 3594 2102 3 FreeSans 24 0 0 0 operand_B[24]
port 92 nsew
flabel metal3 s 3590 2068 3594 2072 3 FreeSans 24 0 0 0 operand_B[25]
port 93 nsew
flabel metal3 s 3590 2298 3594 2302 3 FreeSans 24 0 0 0 operand_B[26]
port 94 nsew
flabel metal3 s 3590 2278 3594 2282 3 FreeSans 24 0 0 0 operand_B[27]
port 95 nsew
flabel metal3 s 3590 2558 3594 2562 3 FreeSans 24 0 0 0 operand_B[28]
port 96 nsew
flabel metal3 s 3590 2708 3594 2712 3 FreeSans 24 0 0 0 operand_B[29]
port 97 nsew
flabel metal3 s 3590 2668 3594 2672 3 FreeSans 24 0 0 0 operand_B[30]
port 98 nsew
flabel metal2 s 3110 3328 3114 3332 3 FreeSans 24 90 0 0 operand_B[31]
port 99 nsew
flabel metal2 s 2662 3328 2666 3332 3 FreeSans 24 90 0 0 operand_B[32]
port 100 nsew
flabel metal2 s 2470 3328 2474 3332 3 FreeSans 24 90 0 0 operand_B[33]
port 101 nsew
flabel metal2 s 2814 3328 2818 3332 3 FreeSans 24 90 0 0 operand_B[34]
port 102 nsew
flabel metal2 s 2926 3328 2930 3332 3 FreeSans 24 90 0 0 operand_B[35]
port 103 nsew
flabel metal2 s 1974 3328 1978 3332 3 FreeSans 24 90 0 0 operand_B[36]
port 104 nsew
flabel metal2 s 2230 3328 2234 3332 3 FreeSans 24 90 0 0 operand_B[37]
port 105 nsew
flabel metal2 s 2278 3328 2282 3332 3 FreeSans 24 90 0 0 operand_B[38]
port 106 nsew
flabel metal2 s 1854 3328 1858 3332 3 FreeSans 24 90 0 0 operand_B[39]
port 107 nsew
flabel metal2 s 1686 3328 1690 3332 3 FreeSans 24 90 0 0 operand_B[40]
port 108 nsew
flabel metal2 s 1550 3328 1554 3332 3 FreeSans 24 90 0 0 operand_B[41]
port 109 nsew
flabel metal2 s 1430 3328 1434 3332 3 FreeSans 24 90 0 0 operand_B[42]
port 110 nsew
flabel metal2 s 1574 3328 1578 3332 3 FreeSans 24 90 0 0 operand_B[43]
port 111 nsew
flabel metal2 s 1726 3328 1730 3332 3 FreeSans 24 90 0 0 operand_B[44]
port 112 nsew
flabel metal2 s 1670 3328 1674 3332 3 FreeSans 24 90 0 0 operand_B[45]
port 113 nsew
flabel metal2 s 1990 3328 1994 3332 3 FreeSans 24 90 0 0 operand_B[46]
port 114 nsew
flabel metal2 s 1646 3328 1650 3332 3 FreeSans 24 90 0 0 operand_B[47]
port 115 nsew
flabel metal2 s 1702 3328 1706 3332 3 FreeSans 24 90 0 0 operand_B[48]
port 116 nsew
flabel metal2 s 1374 3328 1378 3332 3 FreeSans 24 90 0 0 operand_B[49]
port 117 nsew
flabel metal2 s 1286 3328 1290 3332 3 FreeSans 24 90 0 0 operand_B[50]
port 118 nsew
flabel metal2 s 1246 3328 1250 3332 3 FreeSans 24 90 0 0 operand_B[51]
port 119 nsew
flabel metal2 s 734 3328 738 3332 3 FreeSans 24 90 0 0 operand_B[52]
port 120 nsew
flabel metal2 s 646 3328 650 3332 3 FreeSans 24 90 0 0 operand_B[53]
port 121 nsew
flabel metal2 s 750 3328 754 3332 3 FreeSans 24 90 0 0 operand_B[54]
port 122 nsew
flabel metal2 s 670 3328 674 3332 3 FreeSans 24 90 0 0 operand_B[55]
port 123 nsew
flabel metal3 s -26 2648 -22 2652 7 FreeSans 24 0 0 0 operand_B[56]
port 124 nsew
flabel metal3 s -26 2698 -22 2702 7 FreeSans 24 0 0 0 operand_B[57]
port 125 nsew
flabel metal3 s -26 3048 -22 3052 7 FreeSans 24 0 0 0 operand_B[58]
port 126 nsew
flabel metal3 s -26 2868 -22 2872 7 FreeSans 24 0 0 0 operand_B[59]
port 127 nsew
flabel metal3 s -26 2568 -22 2572 7 FreeSans 24 0 0 0 operand_B[60]
port 128 nsew
flabel metal3 s -26 2488 -22 2492 7 FreeSans 24 0 0 0 operand_B[61]
port 129 nsew
flabel metal3 s -26 2548 -22 2552 7 FreeSans 24 0 0 0 operand_B[62]
port 130 nsew
flabel metal2 s 1414 3328 1418 3332 3 FreeSans 24 90 0 0 operand_B[63]
port 131 nsew
flabel metal3 s 3590 1748 3594 1752 3 FreeSans 24 0 0 0 alu_op[0]
port 132 nsew
flabel metal2 s 1142 3328 1146 3332 3 FreeSans 24 90 0 0 alu_op[1]
port 133 nsew
flabel metal3 s 3590 1808 3594 1812 3 FreeSans 24 0 0 0 alu_op[2]
port 134 nsew
flabel metal3 s 3590 1828 3594 1832 3 FreeSans 24 0 0 0 alu_op[3]
port 135 nsew
flabel metal3 s 3590 1548 3594 1552 3 FreeSans 24 0 0 0 result[0]
port 136 nsew
flabel metal3 s 3590 1148 3594 1152 3 FreeSans 24 0 0 0 result[1]
port 137 nsew
flabel metal2 s 2334 -22 2338 -18 7 FreeSans 24 270 0 0 result[2]
port 138 nsew
flabel metal2 s 2366 -22 2370 -18 7 FreeSans 24 270 0 0 result[3]
port 139 nsew
flabel metal2 s 2142 -22 2146 -18 7 FreeSans 24 270 0 0 result[4]
port 140 nsew
flabel metal2 s 2414 -22 2418 -18 7 FreeSans 24 270 0 0 result[5]
port 141 nsew
flabel metal3 s 3590 768 3594 772 3 FreeSans 24 0 0 0 result[6]
port 142 nsew
flabel metal2 s 2766 -22 2770 -18 7 FreeSans 24 270 0 0 result[7]
port 143 nsew
flabel metal3 s 3590 748 3594 752 3 FreeSans 24 0 0 0 result[8]
port 144 nsew
flabel metal3 s 3590 648 3594 652 3 FreeSans 24 0 0 0 result[9]
port 145 nsew
flabel metal3 s 3590 848 3594 852 3 FreeSans 24 0 0 0 result[10]
port 146 nsew
flabel metal3 s 3590 788 3594 792 3 FreeSans 24 0 0 0 result[11]
port 147 nsew
flabel metal3 s 3590 828 3594 832 3 FreeSans 24 0 0 0 result[12]
port 148 nsew
flabel metal3 s 3590 808 3594 812 3 FreeSans 24 0 0 0 result[13]
port 149 nsew
flabel metal3 s 3590 568 3594 572 3 FreeSans 24 0 0 0 result[14]
port 150 nsew
flabel metal3 s 3590 548 3594 552 3 FreeSans 24 0 0 0 result[15]
port 151 nsew
flabel metal3 s 3590 868 3594 872 3 FreeSans 24 0 0 0 result[16]
port 152 nsew
flabel metal3 s 3590 998 3594 1002 3 FreeSans 24 0 0 0 result[17]
port 153 nsew
flabel metal3 s 3590 1168 3594 1172 3 FreeSans 24 0 0 0 result[18]
port 154 nsew
flabel metal3 s 3590 1048 3594 1052 3 FreeSans 24 0 0 0 result[19]
port 155 nsew
flabel metal3 s 3590 3148 3594 3152 3 FreeSans 24 0 0 0 result[20]
port 156 nsew
flabel metal3 s 3590 48 3594 52 3 FreeSans 24 270 0 0 result[21]
port 157 nsew
flabel metal3 s 3590 1848 3594 1852 3 FreeSans 24 0 0 0 result[22]
port 158 nsew
flabel metal3 s 3590 1968 3594 1972 3 FreeSans 24 0 0 0 result[23]
port 159 nsew
flabel metal3 s 3590 1948 3594 1952 3 FreeSans 24 0 0 0 result[24]
port 160 nsew
flabel metal3 s 3590 2048 3594 2052 3 FreeSans 24 0 0 0 result[25]
port 161 nsew
flabel metal3 s 3590 2578 3594 2582 3 FreeSans 24 0 0 0 result[26]
port 162 nsew
flabel metal3 s 3590 2348 3594 2352 3 FreeSans 24 0 0 0 result[27]
port 163 nsew
flabel metal2 s 3542 3328 3546 3332 3 FreeSans 24 90 0 0 result[28]
port 164 nsew
flabel metal2 s 3502 3328 3506 3332 3 FreeSans 24 90 0 0 result[29]
port 165 nsew
flabel metal2 s 3350 3328 3354 3332 3 FreeSans 24 90 0 0 result[30]
port 166 nsew
flabel metal2 s 3326 3328 3330 3332 3 FreeSans 24 90 0 0 result[31]
port 167 nsew
flabel metal2 s 2958 3328 2962 3332 3 FreeSans 24 90 0 0 result[32]
port 168 nsew
flabel metal2 s 2974 3328 2978 3332 3 FreeSans 24 90 0 0 result[33]
port 169 nsew
flabel metal2 s 3230 3328 3234 3332 3 FreeSans 24 90 0 0 result[34]
port 170 nsew
flabel metal2 s 3206 3328 3210 3332 3 FreeSans 24 90 0 0 result[35]
port 171 nsew
flabel metal2 s 3182 3328 3186 3332 3 FreeSans 24 90 0 0 result[36]
port 172 nsew
flabel metal2 s 3158 3328 3162 3332 3 FreeSans 24 90 0 0 result[37]
port 173 nsew
flabel metal2 s 2990 3328 2994 3332 3 FreeSans 24 90 0 0 result[38]
port 174 nsew
flabel metal2 s 3062 3328 3066 3332 3 FreeSans 24 90 0 0 result[39]
port 175 nsew
flabel metal2 s 3014 3328 3018 3332 3 FreeSans 24 90 0 0 result[40]
port 176 nsew
flabel metal2 s 2646 3328 2650 3332 3 FreeSans 24 90 0 0 result[41]
port 177 nsew
flabel metal2 s 2414 3328 2418 3332 3 FreeSans 24 90 0 0 result[42]
port 178 nsew
flabel metal2 s 2502 3328 2506 3332 3 FreeSans 24 90 0 0 result[43]
port 179 nsew
flabel metal2 s 2766 3328 2770 3332 3 FreeSans 24 90 0 0 result[44]
port 180 nsew
flabel metal2 s 2678 3328 2682 3332 3 FreeSans 24 90 0 0 result[45]
port 181 nsew
flabel metal2 s 2598 3328 2602 3332 3 FreeSans 24 90 0 0 result[46]
port 182 nsew
flabel metal2 s 2574 3328 2578 3332 3 FreeSans 24 90 0 0 result[47]
port 183 nsew
flabel metal2 s 2486 3328 2490 3332 3 FreeSans 24 90 0 0 result[48]
port 184 nsew
flabel metal2 s 2342 3328 2346 3332 3 FreeSans 24 90 0 0 result[49]
port 185 nsew
flabel metal2 s 2294 3328 2298 3332 3 FreeSans 24 90 0 0 result[50]
port 186 nsew
flabel metal2 s 2166 3328 2170 3332 3 FreeSans 24 90 0 0 result[51]
port 187 nsew
flabel metal2 s 2094 3328 2098 3332 3 FreeSans 24 90 0 0 result[52]
port 188 nsew
flabel metal2 s 2046 3328 2050 3332 3 FreeSans 24 90 0 0 result[53]
port 189 nsew
flabel metal2 s 526 3328 530 3332 3 FreeSans 24 90 0 0 result[54]
port 190 nsew
flabel metal2 s 2326 3328 2330 3332 3 FreeSans 24 90 0 0 result[55]
port 191 nsew
flabel metal2 s 2310 3328 2314 3332 3 FreeSans 24 90 0 0 result[56]
port 192 nsew
flabel metal2 s 502 3328 506 3332 3 FreeSans 24 90 0 0 result[57]
port 193 nsew
flabel metal2 s 190 3328 194 3332 3 FreeSans 24 90 0 0 result[58]
port 194 nsew
flabel metal3 s -26 3248 -22 3252 7 FreeSans 24 90 0 0 result[59]
port 195 nsew
flabel metal2 s 406 3328 410 3332 3 FreeSans 24 90 0 0 result[60]
port 196 nsew
flabel metal2 s 334 3328 338 3332 3 FreeSans 24 90 0 0 result[61]
port 197 nsew
flabel metal2 s 2438 3328 2442 3332 3 FreeSans 24 90 0 0 result[62]
port 198 nsew
flabel metal2 s 2558 3328 2562 3332 3 FreeSans 24 90 0 0 result[63]
port 199 nsew
flabel metal3 s 3590 2748 3594 2752 3 FreeSans 24 0 0 0 zero_flag
port 200 nsew
flabel metal2 s 174 -22 178 -18 7 FreeSans 24 270 0 0 carry_flag
port 201 nsew
flabel metal2 s 198 -22 202 -18 7 FreeSans 24 270 0 0 overflow_flag
port 202 nsew
<< end >>
