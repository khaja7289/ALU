* NGSPICE file created from ALU_64bit.ext - technology: scmos

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for MUX2X1 abstract view
.subckt MUX2X1 A B S gnd Y vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for OAI22X1 abstract view
.subckt OAI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX2 abstract view
.subckt INVX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX4 abstract view
.subckt BUFX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for XNOR2X1 abstract view
.subckt XNOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX8 abstract view
.subckt INVX8 A gnd Y vdd
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 A gnd Y vdd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for XOR2X1 abstract view
.subckt XOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for DFFPOSX1 abstract view
.subckt DFFPOSX1 Q CLK D gnd vdd
.ends

* Black-box entry subcircuit for INVX4 abstract view
.subckt INVX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for DFFSR abstract view
.subckt DFFSR Q CLK R S D gnd vdd
.ends

.subckt ALU_64bit vdd gnd clk reset operand_A[0] operand_A[1] operand_A[2] operand_A[3]
+ operand_A[4] operand_A[5] operand_A[6] operand_A[7] operand_A[8] operand_A[9] operand_A[10]
+ operand_A[11] operand_A[12] operand_A[13] operand_A[14] operand_A[15] operand_A[16]
+ operand_A[17] operand_A[18] operand_A[19] operand_A[20] operand_A[21] operand_A[22]
+ operand_A[23] operand_A[24] operand_A[25] operand_A[26] operand_A[27] operand_A[28]
+ operand_A[29] operand_A[30] operand_A[31] operand_A[32] operand_A[33] operand_A[34]
+ operand_A[35] operand_A[36] operand_A[37] operand_A[38] operand_A[39] operand_A[40]
+ operand_A[41] operand_A[42] operand_A[43] operand_A[44] operand_A[45] operand_A[46]
+ operand_A[47] operand_A[48] operand_A[49] operand_A[50] operand_A[51] operand_A[52]
+ operand_A[53] operand_A[54] operand_A[55] operand_A[56] operand_A[57] operand_A[58]
+ operand_A[59] operand_A[60] operand_A[61] operand_A[62] operand_A[63] operand_B[0]
+ operand_B[1] operand_B[2] operand_B[3] operand_B[4] operand_B[5] operand_B[6] operand_B[7]
+ operand_B[8] operand_B[9] operand_B[10] operand_B[11] operand_B[12] operand_B[13]
+ operand_B[14] operand_B[15] operand_B[16] operand_B[17] operand_B[18] operand_B[19]
+ operand_B[20] operand_B[21] operand_B[22] operand_B[23] operand_B[24] operand_B[25]
+ operand_B[26] operand_B[27] operand_B[28] operand_B[29] operand_B[30] operand_B[31]
+ operand_B[32] operand_B[33] operand_B[34] operand_B[35] operand_B[36] operand_B[37]
+ operand_B[38] operand_B[39] operand_B[40] operand_B[41] operand_B[42] operand_B[43]
+ operand_B[44] operand_B[45] operand_B[46] operand_B[47] operand_B[48] operand_B[49]
+ operand_B[50] operand_B[51] operand_B[52] operand_B[53] operand_B[54] operand_B[55]
+ operand_B[56] operand_B[57] operand_B[58] operand_B[59] operand_B[60] operand_B[61]
+ operand_B[62] operand_B[63] alu_op[0] alu_op[1] alu_op[2] alu_op[3] result[0] result[1]
+ result[2] result[3] result[4] result[5] result[6] result[7] result[8] result[9]
+ result[10] result[11] result[12] result[13] result[14] result[15] result[16] result[17]
+ result[18] result[19] result[20] result[21] result[22] result[23] result[24] result[25]
+ result[26] result[27] result[28] result[29] result[30] result[31] result[32] result[33]
+ result[34] result[35] result[36] result[37] result[38] result[39] result[40] result[41]
+ result[42] result[43] result[44] result[45] result[46] result[47] result[48] result[49]
+ result[50] result[51] result[52] result[53] result[54] result[55] result[56] result[57]
+ result[58] result[59] result[60] result[61] result[62] result[63] zero_flag carry_flag
+ overflow_flag
XNAND2X1_580 BUFX4_136/Y MUX2X1_110/A gnd OAI21X1_721/C vdd NAND2X1
XNAND2X1_591 BUFX4_191/Y OAI21X1_708/B gnd OAI21X1_736/C vdd NAND2X1
XFILL_17_5_0 gnd vdd FILL
XOAI21X1_360 operand_A[39] INVX2_70/Y NOR2X1_173/Y gnd OAI21X1_361/C vdd OAI21X1
XAND2X2_5 operand_A[30] operand_B[30] gnd AND2X2_5/Y vdd AND2X2
XOAI21X1_382 INVX2_54/Y MUX2X1_3/S OAI21X1_382/C gnd INVX1_164/A vdd OAI21X1
XOAI21X1_371 INVX2_47/Y MUX2X1_7/S OAI21X1_371/C gnd OAI21X1_401/B vdd OAI21X1
XOAI21X1_393 INVX1_169/A OAI21X1_393/B OAI21X1_393/C gnd OAI21X1_393/Y vdd OAI21X1
XFILL_32_3_0 gnd vdd FILL
XAOI21X1_406 BUFX4_79/Y MUX2X1_128/Y INVX8_9/Y gnd OAI22X1_37/C vdd AOI21X1
XFILL_23_3_0 gnd vdd FILL
XMUX2X1_17 operand_A[40] operand_A[39] MUX2X1_6/S gnd MUX2X1_17/Y vdd MUX2X1
XMUX2X1_39 MUX2X1_39/A MUX2X1_39/B BUFX4_22/Y gnd MUX2X1_39/Y vdd MUX2X1
XMUX2X1_28 MUX2X1_28/A MUX2X1_28/B NOR2X1_83/A gnd MUX2X1_28/Y vdd MUX2X1
XFILL_6_4_0 gnd vdd FILL
XFILL_14_3_0 gnd vdd FILL
XINVX1_232 INVX1_232/A gnd INVX1_232/Y vdd INVX1
XINVX1_243 INVX1_243/A gnd INVX1_243/Y vdd INVX1
XINVX1_210 INVX1_210/A gnd INVX1_210/Y vdd INVX1
XINVX1_221 INVX1_221/A gnd INVX1_221/Y vdd INVX1
XOAI21X1_190 MUX2X1_1/Y BUFX4_74/Y OAI21X1_190/C gnd INVX1_90/A vdd OAI21X1
XINVX1_276 BUFX2_26/A gnd INVX1_276/Y vdd INVX1
XINVX1_254 INVX1_254/A gnd INVX1_254/Y vdd INVX1
XNAND2X1_43 INVX2_15/Y INVX1_15/Y gnd NAND2X1_43/Y vdd NAND2X1
XINVX1_298 INVX1_298/A gnd INVX1_298/Y vdd INVX1
XNAND2X1_21 operand_A[6] INVX1_14/Y gnd NAND2X1_23/A vdd NAND2X1
XNAND2X1_32 operand_B[14] INVX2_16/Y gnd INVX2_19/A vdd NAND2X1
XINVX1_287 INVX1_287/A gnd INVX1_287/Y vdd INVX1
XINVX1_265 BUFX2_11/A gnd INVX1_265/Y vdd INVX1
XNAND2X1_10 operand_B[18] INVX4_5/Y gnd NAND2X1_11/B vdd NAND2X1
XNAND2X1_54 operand_B[25] INVX4_8/Y gnd NAND2X1_55/B vdd NAND2X1
XNAND2X1_65 operand_B[23] INVX2_8/Y gnd NAND2X1_65/Y vdd NAND2X1
XNAND2X1_98 BUFX4_120/Y OAI21X1_48/Y gnd OAI21X1_49/C vdd NAND2X1
XNAND2X1_76 XNOR2X1_6/Y XNOR2X1_7/Y gnd NOR2X1_60/A vdd NAND2X1
XNAND2X1_87 BUFX4_67/Y INVX1_91/A gnd OAI21X1_38/C vdd NAND2X1
XAOI21X1_214 AOI21X1_214/A OR2X2_33/Y NAND2X1_485/Y gnd AOI21X1_215/B vdd AOI21X1
XAOI21X1_258 INVX4_24/Y NOR2X1_357/Y BUFX4_30/Y gnd OAI21X1_608/C vdd AOI21X1
XAOI22X1_30 AOI22X1_30/A OAI22X1_26/Y AOI22X1_30/C NOR2X1_281/Y gnd AOI22X1_30/Y vdd
+ AOI22X1
XAOI21X1_247 NOR2X1_345/Y INVX1_246/Y OAI21X1_596/Y gnd OAI21X1_597/C vdd AOI21X1
XAOI21X1_225 INVX1_233/A OAI21X1_500/Y INVX1_236/Y gnd OAI21X1_610/A vdd AOI21X1
XAOI21X1_269 BUFX4_56/Y INVX1_259/A OAI22X1_22/Y gnd NAND2X1_523/B vdd AOI21X1
XAOI21X1_236 INVX8_7/A MUX2X1_57/Y OAI22X1_36/A gnd OAI21X1_588/A vdd AOI21X1
XAOI21X1_203 INVX4_11/Y NAND2X1_477/Y BUFX4_9/Y gnd OAI22X1_32/A vdd AOI21X1
XAOI22X1_41 BUFX4_60/Y XOR2X1_6/Y NAND2X1_42/Y BUFX4_1/Y gnd AOI22X1_41/Y vdd AOI22X1
XAOI22X1_52 BUFX4_148/Y OR2X2_49/B BUFX4_3/Y AOI22X1_52/D gnd AOI22X1_52/Y vdd AOI22X1
XOAI22X1_3 OAI22X1_9/A OR2X2_9/B OAI22X1_3/C OAI22X1_3/D gnd OAI22X1_3/Y vdd OAI22X1
XNAND2X1_409 INVX1_182/A NAND2X1_409/B gnd INVX4_21/A vdd NAND2X1
XNOR2X1_420 NOR2X1_420/A NOR2X1_420/B gnd NOR2X1_421/B vdd NOR2X1
XNOR2X1_431 BUFX4_172/Y INVX1_111/Y gnd NOR2X1_431/Y vdd NOR2X1
XNOR2X1_497 INVX8_7/Y NOR2X1_497/B gnd OAI22X1_33/D vdd NOR2X1
XNOR2X1_442 BUFX4_162/Y NOR2X1_442/B gnd NOR2X1_442/Y vdd NOR2X1
XNOR2X1_453 NOR2X1_453/A NOR2X1_453/B gnd NOR2X1_453/Y vdd NOR2X1
XNOR2X1_464 BUFX4_38/Y NOR2X1_464/B gnd NOR2X1_464/Y vdd NOR2X1
XNOR2X1_475 BUFX4_7/Y NOR2X1_475/B gnd NOR2X1_475/Y vdd NOR2X1
XNOR2X1_486 INVX1_316/Y NOR2X1_486/B gnd NOR2X1_486/Y vdd NOR2X1
XOAI21X1_937 INVX1_326/Y AND2X2_74/A NOR2X1_504/Y gnd OAI21X1_937/Y vdd OAI21X1
XOAI21X1_948 BUFX4_63/Y INVX1_329/Y OAI21X1_948/C gnd NOR2X1_510/B vdd OAI21X1
XOAI21X1_915 OAI21X1_915/A NAND2X1_59/A INVX8_6/A gnd OAI21X1_915/Y vdd OAI21X1
XFILL_20_1_0 gnd vdd FILL
XOAI21X1_926 OAI21X1_926/A BUFX4_169/Y BUFX4_116/Y gnd OAI22X1_36/B vdd OAI21X1
XOAI21X1_904 OAI21X1_904/A NOR2X1_496/Y OR2X2_48/A gnd OAI21X1_905/C vdd OAI21X1
XINVX2_67 operand_B[38] gnd INVX2_67/Y vdd INVX2
XINVX2_78 INVX2_78/A gnd INVX2_78/Y vdd INVX2
XINVX2_56 operand_A[33] gnd INVX2_56/Y vdd INVX2
XINVX2_45 operand_A[32] gnd INVX2_45/Y vdd INVX2
XINVX2_34 INVX2_34/A gnd INVX2_34/Y vdd INVX2
XINVX2_23 operand_B[10] gnd INVX2_23/Y vdd INVX2
XINVX2_12 operand_A[2] gnd INVX2_12/Y vdd INVX2
XFILL_28_2_0 gnd vdd FILL
XINVX2_89 OR2X2_38/A gnd INVX2_89/Y vdd INVX2
XFILL_3_2_0 gnd vdd FILL
XOAI21X1_19 AOI21X1_9/Y OR2X2_1/Y OAI21X1_19/C gnd INVX1_315/A vdd OAI21X1
XFILL_11_1_0 gnd vdd FILL
XFILL_19_2_0 gnd vdd FILL
XNAND2X1_206 INVX4_1/A OAI21X1_94/C gnd NOR2X1_121/B vdd NAND2X1
XNAND2X1_217 MUX2X1_30/S OAI21X1_183/Y gnd OAI21X1_184/C vdd NAND2X1
XNAND2X1_239 BUFX4_133/Y MUX2X1_35/A gnd OAI21X1_209/C vdd NAND2X1
XNAND2X1_228 BUFX4_67/Y INVX1_39/A gnd OAI21X1_195/C vdd NAND2X1
XBUFX4_190 operand_B[1] gnd BUFX4_190/Y vdd BUFX4
XNOR2X1_272 INVX4_23/Y NOR2X1_272/B gnd NOR2X1_273/B vdd NOR2X1
XNOR2X1_261 operand_A[50] operand_B[50] gnd OAI22X1_9/D vdd NOR2X1
XNOR2X1_283 INVX2_53/Y INVX1_218/Y gnd INVX1_222/A vdd NOR2X1
XNOR2X1_250 operand_A[47] INVX1_191/Y gnd NOR2X1_250/Y vdd NOR2X1
XNOR2X1_294 INVX8_7/Y NOR2X1_294/B gnd OAI22X1_32/D vdd NOR2X1
XOAI21X1_701 BUFX4_190/Y operand_A[1] BUFX4_2/Y gnd OAI21X1_702/C vdd OAI21X1
XOAI21X1_712 MUX2X1_95/Y MUX2X1_34/S AND2X2_11/B gnd OAI21X1_714/B vdd OAI21X1
XOAI21X1_723 BUFX4_76/Y MUX2X1_72/Y OAI21X1_723/C gnd INVX1_292/A vdd OAI21X1
XOAI21X1_734 NOR2X1_83/A OAI21X1_734/B OAI21X1_734/C gnd OR2X2_39/A vdd OAI21X1
XOAI21X1_756 BUFX4_162/Y INVX4_7/Y INVX1_297/A gnd INVX1_298/A vdd OAI21X1
XOAI21X1_778 INVX1_297/Y OAI21X1_13/C INVX1_301/Y gnd OAI21X1_781/A vdd OAI21X1
XOAI21X1_745 BUFX4_154/Y NOR2X1_16/Y OAI22X1_7/C gnd OAI21X1_746/C vdd OAI21X1
XOAI21X1_767 BUFX4_97/Y INVX1_266/Y OAI21X1_767/C gnd DFFPOSX1_6/D vdd OAI21X1
XOAI21X1_789 OR2X2_16/A BUFX4_77/Y OAI21X1_789/C gnd OAI21X1_789/Y vdd OAI21X1
XBUFX4_30 INVX8_6/Y gnd BUFX4_30/Y vdd BUFX4
XBUFX4_63 INVX8_17/Y gnd BUFX4_63/Y vdd BUFX4
XBUFX4_52 operand_B[0] gnd MUX2X1_7/S vdd BUFX4
XBUFX4_74 INVX8_1/Y gnd BUFX4_74/Y vdd BUFX4
XBUFX4_41 operand_B[3] gnd BUFX4_41/Y vdd BUFX4
XBUFX4_85 BUFX4_87/A gnd BUFX4_85/Y vdd BUFX4
XBUFX4_96 INVX8_11/Y gnd BUFX4_96/Y vdd BUFX4
XOR2X2_33 OR2X2_33/A OR2X2_33/B gnd OR2X2_33/Y vdd OR2X2
XOR2X2_11 operand_A[37] operand_B[37] gnd OR2X2_11/Y vdd OR2X2
XOR2X2_4 OR2X2_4/A OR2X2_8/B gnd OR2X2_4/Y vdd OR2X2
XOR2X2_44 OR2X2_44/A OR2X2_44/B gnd OR2X2_44/Y vdd OR2X2
XOR2X2_22 OR2X2_22/A OR2X2_39/B gnd OR2X2_22/Y vdd OR2X2
XXNOR2X1_6 operand_A[11] operand_B[11] gnd XNOR2X1_6/Y vdd XNOR2X1
XFILL_26_5_1 gnd vdd FILL
XFILL_25_0_0 gnd vdd FILL
XFILL_1_5_1 gnd vdd FILL
XFILL_0_0_0 gnd vdd FILL
XOAI21X1_531 INVX1_219/Y NOR2X1_286/Y OAI21X1_531/C gnd OAI21X1_531/Y vdd OAI21X1
XOAI21X1_553 INVX1_225/A INVX1_224/A INVX1_226/Y gnd OR2X2_33/A vdd OAI21X1
XOAI21X1_520 INVX1_212/A OAI21X1_520/B AOI22X1_30/A gnd OAI21X1_520/Y vdd OAI21X1
XOAI21X1_564 INVX2_81/A INVX1_232/Y NOR2X1_309/Y gnd OAI21X1_564/Y vdd OAI21X1
XOAI21X1_542 BUFX4_64/Y INVX1_222/Y AOI22X1_22/Y gnd NOR2X1_288/B vdd OAI21X1
XOAI21X1_575 OAI21X1_610/A INVX1_237/Y OAI21X1_584/C gnd NOR2X1_325/B vdd OAI21X1
XINVX8_11 INVX8_11/A gnd INVX8_11/Y vdd INVX8
XINVX1_6 operand_B[16] gnd INVX1_6/Y vdd INVX1
XOAI21X1_597 INVX1_232/A INVX1_247/A OAI21X1_597/C gnd OAI21X1_600/B vdd OAI21X1
XOAI21X1_586 INVX4_9/Y BUFX4_50/Y OAI21X1_64/C gnd MUX2X1_59/B vdd OAI21X1
XNAND2X1_570 BUFX4_72/Y OAI21X1_704/Y gnd OAI21X1_705/C vdd NAND2X1
XNAND2X1_581 BUFX4_71/Y INVX1_284/Y gnd OAI21X1_722/C vdd NAND2X1
XNAND2X1_592 BUFX4_125/Y MUX2X1_114/A gnd OAI21X1_737/C vdd NAND2X1
XFILL_8_1_0 gnd vdd FILL
XFILL_17_5_1 gnd vdd FILL
XFILL_16_0_0 gnd vdd FILL
XOAI21X1_361 INVX2_69/Y operand_B[39] OAI21X1_361/C gnd NOR2X1_184/A vdd OAI21X1
XAND2X2_6 AND2X2_6/A INVX1_75/A gnd AND2X2_6/Y vdd AND2X2
XOAI21X1_394 INVX1_162/A AND2X2_16/B OAI21X1_394/C gnd NOR2X1_203/A vdd OAI21X1
XOAI21X1_372 INVX1_159/Y BUFX4_75/Y OAI21X1_372/C gnd OAI21X1_372/Y vdd OAI21X1
XOAI21X1_383 INVX1_164/Y BUFX4_190/Y OAI21X1_383/C gnd INVX1_165/A vdd OAI21X1
XOAI21X1_350 INVX1_121/Y MUX2X1_27/S OAI21X1_350/C gnd INVX1_196/A vdd OAI21X1
XFILL_32_3_1 gnd vdd FILL
XAOI21X1_407 BUFX4_141/Y XNOR2X1_48/Y NAND2X1_649/Y gnd AOI22X1_57/C vdd AOI21X1
XFILL_23_3_1 gnd vdd FILL
XMUX2X1_18 operand_A[44] operand_A[43] MUX2X1_3/S gnd MUX2X1_18/Y vdd MUX2X1
XMUX2X1_29 MUX2X1_29/A MUX2X1_29/B BUFX4_35/Y gnd MUX2X1_29/Y vdd MUX2X1
XFILL_6_4_1 gnd vdd FILL
XFILL_14_3_1 gnd vdd FILL
XINVX1_222 INVX1_222/A gnd INVX1_222/Y vdd INVX1
XINVX1_244 INVX1_244/A gnd INVX1_244/Y vdd INVX1
XINVX1_233 INVX1_233/A gnd INVX1_233/Y vdd INVX1
XINVX1_211 operand_A[51] gnd INVX1_211/Y vdd INVX1
XINVX1_200 INVX1_200/A gnd INVX1_200/Y vdd INVX1
XINVX1_255 INVX1_255/A gnd INVX1_255/Y vdd INVX1
XAOI22X1_1 AOI22X1_1/A AOI22X1_1/B INVX1_32/Y NOR2X1_67/Y gnd AOI22X1_1/Y vdd AOI22X1
XOAI21X1_180 BUFX4_71/Y MUX2X1_9/Y OAI21X1_180/C gnd MUX2X1_24/B vdd OAI21X1
XINVX1_277 BUFX2_25/A gnd INVX1_277/Y vdd INVX1
XOAI21X1_191 INVX1_44/Y BUFX4_76/Y OAI21X1_191/C gnd OAI21X1_290/B vdd OAI21X1
XINVX1_266 BUFX2_8/A gnd INVX1_266/Y vdd INVX1
XNAND2X1_44 operand_B[26] operand_A[26] gnd OAI21X1_20/C vdd NAND2X1
XNAND2X1_55 NAND2X1_55/A NAND2X1_55/B gnd NAND2X1_59/A vdd NAND2X1
XNAND2X1_66 INVX1_28/Y NAND2X1_66/B gnd NAND2X1_66/Y vdd NAND2X1
XNAND2X1_77 INVX2_17/A INVX1_17/A gnd NOR2X1_60/B vdd NAND2X1
XNAND2X1_22 operand_B[6] INVX2_13/Y gnd INVX1_281/A vdd NAND2X1
XINVX1_288 INVX1_288/A gnd INVX1_288/Y vdd INVX1
XNAND2X1_33 INVX2_18/A INVX2_19/A gnd OR2X2_45/B vdd NAND2X1
XINVX1_299 INVX1_299/A gnd INVX1_299/Y vdd INVX1
XNAND2X1_11 NAND2X1_9/Y NAND2X1_11/B gnd OR2X2_47/B vdd NAND2X1
XNAND2X1_88 MUX2X1_1/S operand_A[19] gnd OAI21X1_39/C vdd NAND2X1
XNAND2X1_99 BUFX4_17/Y INVX1_42/Y gnd OAI21X1_50/C vdd NAND2X1
XAOI21X1_215 OAI21X1_552/Y AOI21X1_215/B NOR2X1_302/Y gnd DFFPOSX1_56/D vdd AOI21X1
XAOI21X1_248 OAI21X1_472/C OAI21X1_598/Y INVX1_231/A gnd OAI21X1_599/A vdd AOI21X1
XAOI22X1_20 BUFX4_153/Y NOR2X1_258/B BUFX4_58/Y INVX1_204/A gnd AND2X2_29/A vdd AOI22X1
XAOI21X1_259 INVX2_89/Y OAI21X1_610/Y NAND2X1_516/Y gnd AOI21X1_262/A vdd AOI21X1
XAOI21X1_237 BUFX4_111/Y OAI22X1_36/D OAI21X1_587/Y gnd OAI21X1_588/C vdd AOI21X1
XAOI22X1_53 BUFX4_148/Y NOR2X1_11/Y AOI21X1_4/A BUFX4_3/Y gnd NAND3X1_71/A vdd AOI22X1
XAOI21X1_226 INVX4_11/Y NAND2X1_497/Y BUFX4_9/Y gnd OAI22X1_35/A vdd AOI21X1
XAOI21X1_204 INVX8_7/A OAI21X1_548/Y OAI22X1_32/A gnd OAI21X1_551/A vdd AOI21X1
XAOI22X1_31 BUFX4_12/Y INVX1_269/Y AOI22X1_31/C AOI22X1_31/D gnd DFFPOSX1_1/D vdd
+ AOI22X1
XAOI22X1_42 BUFX4_15/Y INVX1_262/Y AND2X2_60/Y AOI22X1_42/D gnd AOI22X1_42/Y vdd AOI22X1
XOAI22X1_4 OAI22X1_9/A INVX4_19/Y OAI22X1_4/C INVX8_15/Y gnd OAI22X1_4/Y vdd OAI22X1
XNOR2X1_410 XOR2X1_3/Y NOR2X1_410/B gnd AND2X2_46/A vdd NOR2X1
XNOR2X1_421 NOR2X1_421/A NOR2X1_421/B gnd NOR2X1_421/Y vdd NOR2X1
XOAI21X1_916 OAI21X1_34/A NAND2X1_59/B NAND2X1_58/A gnd XNOR2X1_47/A vdd OAI21X1
XNOR2X1_498 OR2X2_48/A BUFX2_27/A gnd NOR2X1_498/Y vdd NOR2X1
XOAI21X1_905 OR2X2_48/A INVX1_277/Y OAI21X1_905/C gnd OAI21X1_905/Y vdd OAI21X1
XNOR2X1_487 BUFX4_7/Y NOR2X1_487/B gnd OAI22X1_29/A vdd NOR2X1
XNOR2X1_432 MUX2X1_23/S NOR2X1_432/B gnd NOR2X1_432/Y vdd NOR2X1
XNOR2X1_476 NOR2X1_40/Y INVX1_313/A gnd NOR2X1_476/Y vdd NOR2X1
XNOR2X1_443 NOR2X1_22/A operand_A[5] gnd INVX1_301/A vdd NOR2X1
XNOR2X1_454 NOR2X1_454/A NOR2X1_454/B gnd AND2X2_58/B vdd NOR2X1
XNOR2X1_465 BUFX4_24/Y NOR2X1_465/B gnd NOR2X1_465/Y vdd NOR2X1
XOAI21X1_949 BUFX4_158/Y NOR2X1_3/A BUFX4_99/Y gnd NOR2X1_510/A vdd OAI21X1
XOAI21X1_938 OAI21X1_34/Y NOR2X1_3/B BUFX4_141/Y gnd OAI21X1_938/Y vdd OAI21X1
XOAI21X1_927 operand_B[26] operand_A[26] BUFX4_6/Y gnd OAI21X1_928/C vdd OAI21X1
XFILL_20_1_1 gnd vdd FILL
XINVX2_68 OR2X2_12/B gnd INVX2_68/Y vdd INVX2
XINVX2_79 INVX2_79/A gnd OR2X2_33/B vdd INVX2
XINVX2_35 operand_A[30] gnd INVX2_35/Y vdd INVX2
XINVX2_46 operand_A[44] gnd INVX2_46/Y vdd INVX2
XINVX2_57 INVX2_57/A gnd INVX2_57/Y vdd INVX2
XINVX2_24 operand_A[9] gnd INVX2_24/Y vdd INVX2
XINVX2_13 operand_A[6] gnd INVX2_13/Y vdd INVX2
XFILL_28_2_1 gnd vdd FILL
XFILL_3_2_1 gnd vdd FILL
XFILL_11_1_1 gnd vdd FILL
XFILL_19_2_1 gnd vdd FILL
XNAND2X1_207 INVX1_33/A NOR2X1_121/Y gnd NOR2X1_122/B vdd NAND2X1
XNAND2X1_218 BUFX4_38/Y INVX1_88/Y gnd OAI21X1_185/C vdd NAND2X1
XNAND2X1_229 BUFX4_119/Y INVX1_128/A gnd OAI21X1_196/C vdd NAND2X1
XNOR2X1_240 BUFX4_102/Y BUFX2_51/A gnd NOR2X1_240/Y vdd NOR2X1
XNOR2X1_251 OR2X2_30/Y NOR2X1_251/B gnd NOR2X1_251/Y vdd NOR2X1
XBUFX4_191 operand_B[1] gnd BUFX4_191/Y vdd BUFX4
XBUFX4_180 operand_B[4] gnd MUX2X1_34/S vdd BUFX4
XNOR2X1_295 BUFX4_98/Y OR2X2_37/A gnd NOR2X1_295/Y vdd NOR2X1
XNOR2X1_273 NOR2X1_273/A NOR2X1_273/B gnd NOR2X1_273/Y vdd NOR2X1
XNOR2X1_284 operand_A[53] operand_B[53] gnd INVX1_223/A vdd NOR2X1
XNOR2X1_262 INVX2_41/Y INVX2_76/Y gnd NOR2X1_273/A vdd NOR2X1
XOAI21X1_735 BUFX4_190/Y MUX2X1_79/Y OAI21X1_735/C gnd INVX1_295/A vdd OAI21X1
XOAI21X1_757 XNOR2X1_20/Y INVX1_298/Y OAI21X1_757/C gnd NAND3X1_61/C vdd OAI21X1
XOAI21X1_713 XOR2X1_3/Y NOR2X1_112/Y OAI21X1_713/C gnd OAI21X1_714/C vdd OAI21X1
XOAI21X1_702 BUFX4_62/Y INVX1_289/Y OAI21X1_702/C gnd OAI21X1_702/Y vdd OAI21X1
XOAI21X1_746 BUFX4_35/Y operand_A[3] OAI21X1_746/C gnd OAI21X1_746/Y vdd OAI21X1
XOAI21X1_724 MUX2X1_27/S MUX2X1_111/A OAI21X1_724/C gnd OAI21X1_727/A vdd OAI21X1
XOAI21X1_779 OAI21X1_781/A XNOR2X1_19/Y BUFX4_105/Y gnd OAI21X1_779/Y vdd OAI21X1
XOAI21X1_768 INVX1_292/Y MUX2X1_27/S OAI21X1_768/C gnd OAI21X1_852/B vdd OAI21X1
XBUFX4_20 INVX8_2/Y gnd BUFX4_20/Y vdd BUFX4
XBUFX4_64 INVX8_17/Y gnd BUFX4_64/Y vdd BUFX4
XBUFX4_75 INVX8_1/Y gnd BUFX4_75/Y vdd BUFX4
XBUFX4_31 INVX8_6/Y gnd BUFX4_31/Y vdd BUFX4
XBUFX4_53 operand_B[0] gnd BUFX4_53/Y vdd BUFX4
XBUFX4_42 operand_B[3] gnd BUFX4_42/Y vdd BUFX4
XBUFX4_86 BUFX4_87/A gnd BUFX4_86/Y vdd BUFX4
XBUFX4_97 DFFSR_1/Q gnd BUFX4_97/Y vdd BUFX4
XFILL_10_1 gnd vdd FILL
XOR2X2_12 OR2X2_12/A OR2X2_12/B gnd OR2X2_12/Y vdd OR2X2
XOR2X2_34 OR2X2_34/A OR2X2_34/B gnd OR2X2_34/Y vdd OR2X2
XOR2X2_23 OR2X2_23/A OR2X2_23/B gnd OR2X2_23/Y vdd OR2X2
XOR2X2_45 OR2X2_45/A OR2X2_45/B gnd OR2X2_45/Y vdd OR2X2
XOR2X2_5 OR2X2_5/A OR2X2_5/B gnd OR2X2_5/Y vdd OR2X2
XXNOR2X1_7 operand_B[10] operand_A[10] gnd XNOR2X1_7/Y vdd XNOR2X1
XFILL_25_0_1 gnd vdd FILL
XINVX8_12 INVX8_12/A gnd BUFX4_9/A vdd INVX8
XFILL_0_0_1 gnd vdd FILL
XOAI21X1_543 INVX1_216/A NOR2X1_307/B OAI21X1_563/A gnd OAI21X1_544/B vdd OAI21X1
XOAI21X1_532 OAI22X1_11/D AND2X2_32/Y OAI21X1_532/C gnd OAI21X1_533/C vdd OAI21X1
XOAI21X1_510 XNOR2X1_37/A INVX4_23/A OAI21X1_520/B gnd XNOR2X1_38/A vdd OAI21X1
XOAI21X1_521 OAI21X1_565/A NOR2X1_311/B NOR2X1_312/B gnd OAI21X1_532/C vdd OAI21X1
XOAI21X1_565 OAI21X1_565/A INVX1_233/Y INVX1_236/A gnd OAI21X1_566/B vdd OAI21X1
XOAI21X1_598 AOI21X1_50/Y AOI21X1_47/C NOR2X1_346/Y gnd OAI21X1_598/Y vdd OAI21X1
XOAI21X1_576 INVX4_13/Y MUX2X1_1/S OAI21X1_576/C gnd INVX1_238/A vdd OAI21X1
XOAI21X1_587 OAI21X1_926/A BUFX4_174/Y AND2X2_42/Y gnd OAI21X1_587/Y vdd OAI21X1
XOAI21X1_554 INVX1_66/Y BUFX4_35/Y OR2X2_43/B gnd OAI21X1_555/C vdd OAI21X1
XINVX1_7 operand_B[19] gnd INVX1_7/Y vdd INVX1
XFILL_8_1_1 gnd vdd FILL
XNAND2X1_560 MUX2X1_7/S operand_A[9] gnd OAI21X1_682/C vdd NAND2X1
XNAND2X1_593 NOR2X1_82/A OAI21X1_710/B gnd OAI21X1_739/C vdd NAND2X1
XNAND2X1_582 BUFX4_76/Y OAI21X1_680/Y gnd OAI21X1_723/C vdd NAND2X1
XNAND2X1_571 BUFX4_38/Y MUX2X1_118/A gnd NAND2X1_571/Y vdd NAND2X1
XFILL_16_0_1 gnd vdd FILL
XOAI21X1_395 AND2X2_17/Y NOR2X1_203/A INVX1_169/Y gnd AND2X2_19/A vdd OAI21X1
XOAI21X1_362 INVX1_126/Y INVX1_157/Y AND2X2_27/A gnd OAI21X1_362/Y vdd OAI21X1
XAND2X2_7 AND2X2_7/A BUFX4_21/Y gnd AND2X2_7/Y vdd AND2X2
XOAI21X1_384 INVX1_165/Y NOR2X1_83/A OAI21X1_384/C gnd MUX2X1_43/B vdd OAI21X1
XOAI21X1_373 INVX1_131/Y MUX2X1_62/S OAI21X1_373/C gnd INVX1_160/A vdd OAI21X1
XOAI21X1_340 INVX1_46/Y BUFX4_23/Y OAI21X1_340/C gnd INVX1_147/A vdd OAI21X1
XOAI21X1_351 INVX1_64/Y BUFX4_23/Y OAI21X1_351/C gnd NOR2X1_300/B vdd OAI21X1
XNAND2X1_390 BUFX4_23/Y INVX1_120/Y gnd OAI21X1_411/C vdd NAND2X1
XAOI21X1_408 NOR2X1_3/B OAI21X1_34/Y OAI21X1_938/Y gnd NOR2X1_506/A vdd AOI21X1
XMUX2X1_19 operand_A[36] operand_A[35] MUX2X1_4/S gnd MUX2X1_19/Y vdd MUX2X1
XAOI22X1_2 BUFX4_148/Y AND2X2_5/Y INVX4_1/Y BUFX4_57/Y gnd NAND3X1_3/B vdd AOI22X1
XINVX1_212 INVX1_212/A gnd INVX1_212/Y vdd INVX1
XINVX1_223 INVX1_223/A gnd INVX1_223/Y vdd INVX1
XINVX1_201 INVX1_201/A gnd INVX1_201/Y vdd INVX1
XINVX1_256 operand_B[62] gnd INVX1_256/Y vdd INVX1
XINVX1_245 operand_B[60] gnd INVX1_245/Y vdd INVX1
XOAI21X1_170 INVX2_29/Y operand_A[27] AOI22X1_1/B gnd OAI21X1_171/C vdd OAI21X1
XOAI21X1_181 BUFX4_72/Y MUX2X1_6/Y OAI21X1_181/C gnd MUX2X1_24/A vdd OAI21X1
XINVX1_234 INVX1_234/A gnd INVX1_234/Y vdd INVX1
XINVX1_278 INVX1_278/A gnd INVX1_278/Y vdd INVX1
XOAI21X1_192 INVX1_90/Y MUX2X1_2/S OAI21X1_192/C gnd OAI21X1_369/A vdd OAI21X1
XINVX1_289 NOR2X1_15/Y gnd INVX1_289/Y vdd INVX1
XINVX1_267 BUFX2_7/A gnd INVX1_267/Y vdd INVX1
XNAND2X1_45 operand_B[27] INVX2_30/Y gnd AOI22X1_1/A vdd NAND2X1
XNAND2X1_56 operand_A[24] INVX1_24/Y gnd NAND2X1_58/A vdd NAND2X1
XNAND2X1_78 NOR2X1_59/Y NOR2X1_60/Y gnd OAI21X1_32/B vdd NAND2X1
XNAND2X1_34 operand_A[13] INVX1_18/Y gnd NAND2X1_36/A vdd NAND2X1
XNAND2X1_23 NAND2X1_23/A INVX1_281/A gnd OAI21X1_10/C vdd NAND2X1
XNAND2X1_67 BUFX4_190/Y INVX2_9/Y gnd INVX1_279/A vdd NAND2X1
XNAND2X1_89 MUX2X1_6/S operand_A[21] gnd OAI21X1_40/C vdd NAND2X1
XNAND2X1_12 XOR2X1_2/Y OR2X2_47/B gnd OAI21X1_3/A vdd NAND2X1
XAOI21X1_216 AND2X2_33/Y INVX1_229/Y AND2X2_35/Y gnd AND2X2_36/B vdd AOI21X1
XAOI21X1_205 BUFX4_149/Y AND2X2_33/Y OAI22X1_13/Y gnd AND2X2_34/A vdd AOI21X1
XAOI21X1_238 BUFX4_143/Y NOR2X1_332/Y OAI21X1_588/Y gnd AOI21X1_239/B vdd AOI21X1
XAOI21X1_249 OAI21X1_597/C OAI21X1_599/Y INVX2_88/Y gnd NOR2X1_357/B vdd AOI21X1
XAOI22X1_21 BUFX4_56/Y INVX1_212/A BUFX4_4/Y INVX1_214/Y gnd NAND3X1_30/B vdd AOI22X1
XAOI22X1_10 BUFX4_153/Y NOR2X1_190/B BUFX4_58/Y INVX1_162/A gnd AOI22X1_10/Y vdd AOI22X1
XAOI22X1_54 BUFX4_13/Y INVX1_276/Y AOI22X1_54/C AOI22X1_54/D gnd AOI22X1_54/Y vdd
+ AOI22X1
XAOI21X1_227 BUFX4_167/Y MUX2X1_55/Y INVX8_7/Y gnd AOI21X1_228/B vdd AOI21X1
XAOI22X1_43 BUFX4_60/Y XNOR2X1_41/B INVX1_21/Y BUFX4_1/Y gnd AOI22X1_43/Y vdd AOI22X1
XAOI22X1_32 BUFX4_12/Y INVX1_268/Y AND2X2_53/Y NOR2X1_429/Y gnd DFFPOSX1_2/D vdd AOI22X1
XOAI22X1_5 BUFX4_61/Y INVX2_63/A OAI22X1_9/C OAI22X1_5/D gnd OAI22X1_5/Y vdd OAI22X1
XNOR2X1_411 INVX1_248/A OR2X2_38/Y gnd NOR2X1_411/Y vdd NOR2X1
XNOR2X1_422 operand_A[46] INVX1_184/Y gnd NOR2X1_422/Y vdd NOR2X1
XNOR2X1_433 NOR2X1_433/A NOR2X1_433/B gnd NOR2X1_433/Y vdd NOR2X1
XNOR2X1_400 NOR2X1_400/A NOR2X1_400/B gnd NOR2X1_400/Y vdd NOR2X1
XOAI21X1_928 BUFX4_63/Y OAI21X1_20/C OAI21X1_928/C gnd NOR2X1_500/B vdd OAI21X1
XNOR2X1_499 NOR2X1_499/A NOR2X1_499/B gnd NOR2X1_499/Y vdd NOR2X1
XOAI21X1_939 OAI21X1_939/A BUFX4_169/Y INVX8_4/A gnd OAI22X1_38/B vdd OAI21X1
XOAI21X1_906 operand_B[22] INVX4_3/Y OAI21X1_906/C gnd OAI21X1_907/B vdd OAI21X1
XOAI21X1_917 OAI21X1_917/A BUFX4_169/Y OR2X2_40/B gnd OAI22X1_35/B vdd OAI21X1
XNOR2X1_477 BUFX4_83/Y OAI22X1_8/B gnd NOR2X1_477/Y vdd NOR2X1
XNOR2X1_455 BUFX4_179/Y NOR2X1_455/B gnd NOR2X1_456/B vdd NOR2X1
XNOR2X1_444 INVX8_15/Y NOR2X1_444/B gnd NOR2X1_444/Y vdd NOR2X1
XNOR2X1_466 NOR2X1_22/A AND2X2_61/Y gnd NOR2X1_466/Y vdd NOR2X1
XNOR2X1_488 NOR2X1_488/A NOR2X1_488/B gnd NOR2X1_488/Y vdd NOR2X1
XINVX2_69 operand_A[39] gnd INVX2_69/Y vdd INVX2
XINVX2_47 operand_A[40] gnd INVX2_47/Y vdd INVX2
XINVX2_36 INVX2_36/A gnd INVX2_36/Y vdd INVX2
XINVX2_25 operand_B[9] gnd INVX2_25/Y vdd INVX2
XINVX2_58 INVX2_58/A gnd INVX2_58/Y vdd INVX2
XINVX2_14 operand_A[5] gnd INVX2_14/Y vdd INVX2
XFILL_30_4_0 gnd vdd FILL
XNAND2X1_208 BUFX4_68/Y OAI21X1_69/B gnd OAI21X1_175/C vdd NAND2X1
XNAND2X1_219 BUFX4_164/Y MUX2X1_123/A gnd OAI21X1_186/C vdd NAND2X1
XNOR2X1_263 OAI22X1_9/D NOR2X1_273/A gnd INVX4_23/A vdd NOR2X1
XNOR2X1_285 INVX1_223/A INVX1_222/A gnd INVX1_219/A vdd NOR2X1
XNOR2X1_241 operand_A[48] operand_B[48] gnd INVX1_202/A vdd NOR2X1
XNOR2X1_230 operand_A[46] operand_B[46] gnd NOR2X1_231/A vdd NOR2X1
XBUFX4_170 INVX8_10/Y gnd NOR2X1_87/B vdd BUFX4
XNOR2X1_252 NOR2X1_87/B NOR2X1_252/B gnd NOR2X1_253/A vdd NOR2X1
XBUFX4_192 operand_B[1] gnd BUFX4_192/Y vdd BUFX4
XBUFX4_181 operand_B[4] gnd OR2X2_7/B vdd BUFX4
XNOR2X1_274 INVX8_7/Y MUX2X1_46/Y gnd NOR2X1_274/Y vdd NOR2X1
XNOR2X1_296 operand_A[55] operand_B[55] gnd INVX1_229/A vdd NOR2X1
XFILL_21_4_0 gnd vdd FILL
XOAI21X1_703 BUFX4_72/Y OAI21X1_703/B OAI21X1_703/C gnd OAI21X1_703/Y vdd OAI21X1
XOAI21X1_725 BUFX4_72/Y MUX2X1_69/A OAI21X1_725/C gnd MUX2X1_111/B vdd OAI21X1
XOAI21X1_758 AOI21X1_51/Y INVX2_92/Y NAND2X1_26/A gnd OAI21X1_759/B vdd OAI21X1
XOAI21X1_747 BUFX4_134/Y MUX2X1_76/Y OAI21X1_747/C gnd OAI21X1_747/Y vdd OAI21X1
XOAI21X1_769 BUFX4_38/Y MUX2X1_110/Y OAI21X1_769/C gnd OAI21X1_770/B vdd OAI21X1
XOAI21X1_714 OAI21X1_714/A OAI21X1_714/B OAI21X1_714/C gnd NOR2X1_429/B vdd OAI21X1
XOAI21X1_736 BUFX4_192/Y MUX2X1_80/Y OAI21X1_736/C gnd MUX2X1_114/A vdd OAI21X1
XFILL_29_5_0 gnd vdd FILL
XFILL_4_5_0 gnd vdd FILL
XFILL_12_4_0 gnd vdd FILL
XINVX8_1 INVX8_1/A gnd INVX8_1/Y vdd INVX8
XBUFX4_32 INVX8_6/Y gnd BUFX4_32/Y vdd BUFX4
XBUFX4_10 BUFX4_9/A gnd BUFX4_10/Y vdd BUFX4
XBUFX4_21 INVX8_2/Y gnd BUFX4_21/Y vdd BUFX4
XBUFX4_43 operand_B[0] gnd BUFX4_43/Y vdd BUFX4
XBUFX4_98 DFFSR_1/Q gnd BUFX4_98/Y vdd BUFX4
XBUFX4_65 INVX8_17/Y gnd BUFX4_65/Y vdd BUFX4
XBUFX4_54 operand_B[0] gnd MUX2X1_3/S vdd BUFX4
XBUFX4_76 INVX8_1/Y gnd BUFX4_76/Y vdd BUFX4
XBUFX4_87 BUFX4_87/A gnd INVX8_15/A vdd BUFX4
XOR2X2_6 operand_A[33] operand_B[33] gnd OR2X2_6/Y vdd OR2X2
XOR2X2_24 OR2X2_24/A OR2X2_24/B gnd OR2X2_24/Y vdd OR2X2
XOR2X2_35 OR2X2_35/A OR2X2_8/B gnd OR2X2_35/Y vdd OR2X2
XOR2X2_13 OR2X2_13/A OR2X2_13/B gnd OR2X2_13/Y vdd OR2X2
XXNOR2X1_8 operand_A[9] operand_B[9] gnd INVX2_17/A vdd XNOR2X1
XOR2X2_46 OR2X2_46/A OR2X2_46/B gnd OR2X2_46/Y vdd OR2X2
XINVX8_13 OR2X2_8/B gnd INVX8_13/Y vdd INVX8
XOAI21X1_544 INVX1_224/A OAI21X1_544/B OAI21X1_544/C gnd OAI21X1_544/Y vdd OAI21X1
XOAI21X1_522 INVX2_78/Y OAI21X1_532/C OAI21X1_522/C gnd NAND3X1_31/A vdd OAI21X1
XOAI21X1_533 INVX2_40/Y operand_B[52] OAI21X1_533/C gnd XNOR2X1_39/A vdd OAI21X1
XOAI21X1_599 OAI21X1_599/A OAI21X1_599/B INVX1_247/Y gnd OAI21X1_599/Y vdd OAI21X1
XOAI21X1_566 INVX2_81/Y OAI21X1_566/B OAI21X1_566/C gnd AND2X2_38/A vdd OAI21X1
XOAI21X1_500 AOI21X1_62/B INVX1_199/A OAI21X1_500/C gnd OAI21X1_500/Y vdd OAI21X1
XOAI21X1_511 INVX1_211/Y MUX2X1_3/S OAI21X1_511/C gnd OAI21X1_511/Y vdd OAI21X1
XOAI21X1_577 BUFX4_70/Y OAI21X1_577/B OAI21X1_577/C gnd MUX2X1_62/B vdd OAI21X1
XOAI21X1_588 OAI21X1_588/A BUFX4_112/Y OAI21X1_588/C gnd OAI21X1_588/Y vdd OAI21X1
XINVX1_8 operand_B[23] gnd INVX1_8/Y vdd INVX1
XOAI21X1_555 INVX1_150/A BUFX4_179/Y OAI21X1_555/C gnd NOR2X1_497/B vdd OAI21X1
XNAND2X1_550 operand_B[32] INVX2_45/Y gnd OAI21X1_666/B vdd NAND2X1
XNAND2X1_561 MUX2X1_23/S OAI21X1_683/Y gnd OAI21X1_684/C vdd NAND2X1
XNAND2X1_572 BUFX4_191/Y MUX2X1_79/Y gnd OAI21X1_708/C vdd NAND2X1
XNAND2X1_594 NAND2X1_594/A OAI21X1_746/Y gnd NOR2X1_437/A vdd NAND2X1
XNAND2X1_583 BUFX4_125/Y INVX1_292/Y gnd OAI21X1_724/C vdd NAND2X1
XFILL_9_1 gnd vdd FILL
XFILL_26_3_0 gnd vdd FILL
XFILL_1_3_0 gnd vdd FILL
XOAI21X1_330 OAI22X1_5/D INVX2_63/Y INVX2_65/A gnd NOR2X1_420/A vdd OAI21X1
XOAI21X1_341 INVX1_147/Y MUX2X1_25/S OAI21X1_341/C gnd OAI22X1_6/C vdd OAI21X1
XOAI21X1_363 INVX1_154/A INVX1_163/A OAI21X1_363/C gnd OAI21X1_364/C vdd OAI21X1
XAND2X2_8 AND2X2_8/A INVX8_13/Y gnd AND2X2_8/Y vdd AND2X2
XOAI21X1_374 BUFX4_18/Y OAI21X1_374/B OAI21X1_374/C gnd NOR2X1_316/B vdd OAI21X1
XOAI21X1_352 INVX1_149/Y BUFX4_20/Y OAI21X1_352/C gnd INVX1_150/A vdd OAI21X1
XOAI21X1_396 MUX2X1_2/B BUFX4_131/Y BUFX4_42/Y gnd OAI21X1_397/C vdd OAI21X1
XOAI21X1_385 BUFX4_37/Y MUX2X1_26/B OAI21X1_385/C gnd OAI22X1_15/B vdd OAI21X1
XNAND2X1_391 BUFX4_69/Y OAI21X1_412/Y gnd OAI21X1_413/C vdd NAND2X1
XNAND2X1_380 BUFX4_36/Y OAI21X1_213/B gnd OAI21X1_385/C vdd NAND2X1
XFILL_9_4_0 gnd vdd FILL
XFILL_17_3_0 gnd vdd FILL
XAOI21X1_409 BUFX4_80/Y MUX2X1_129/Y INVX8_9/Y gnd OAI22X1_38/D vdd AOI21X1
XAOI22X1_3 BUFX4_148/Y INVX1_75/Y BUFX4_6/Y AND2X2_6/A gnd AOI22X1_3/Y vdd AOI22X1
XOAI21X1_171 INVX1_32/A NOR2X1_70/A OAI21X1_171/C gnd AOI21X1_60/A vdd OAI21X1
XOAI21X1_182 INVX1_87/Y BUFX4_71/Y OAI21X1_182/C gnd OAI21X1_299/B vdd OAI21X1
XOAI21X1_160 AOI21X1_51/Y OR2X2_3/Y AOI21X1_52/Y gnd AOI21X1_55/B vdd OAI21X1
XINVX1_224 INVX1_224/A gnd INVX1_224/Y vdd INVX1
XINVX1_202 INVX1_202/A gnd INVX1_202/Y vdd INVX1
XINVX1_246 INVX1_246/A gnd INVX1_246/Y vdd INVX1
XINVX1_257 INVX1_257/A gnd INVX1_257/Y vdd INVX1
XINVX1_235 operand_B[57] gnd INVX1_235/Y vdd INVX1
XINVX1_213 INVX1_213/A gnd INVX1_213/Y vdd INVX1
XINVX1_279 INVX1_279/A gnd INVX1_279/Y vdd INVX1
XOAI21X1_193 BUFX4_41/Y OAI21X1_375/B OAI21X1_193/C gnd MUX2X1_25/B vdd OAI21X1
XINVX1_268 BUFX2_4/A gnd INVX1_268/Y vdd INVX1
XNAND2X1_46 operand_A[27] INVX2_29/Y gnd NAND2X1_47/B vdd NAND2X1
XNAND2X1_57 operand_B[24] INVX2_32/Y gnd NAND2X1_58/B vdd NAND2X1
XNAND2X1_79 operand_B[9] INVX2_24/Y gnd NAND2X1_79/Y vdd NAND2X1
XNAND2X1_35 operand_B[13] INVX2_20/Y gnd NAND2X1_36/B vdd NAND2X1
XNAND2X1_68 MUX2X1_4/S INVX1_29/Y gnd NAND2X1_68/Y vdd NAND2X1
XNAND2X1_24 operand_A[4] BUFX4_162/Y gnd NAND2X1_26/A vdd NAND2X1
XNAND2X1_13 INVX1_5/Y INVX4_6/Y gnd AOI21X1_2/A vdd NAND2X1
XFILL_32_1_0 gnd vdd FILL
XAOI21X1_239 OAI21X1_583/Y AOI21X1_239/B NOR2X1_335/Y gnd DFFPOSX1_59/D vdd AOI21X1
XAOI21X1_217 INVX1_231/Y AND2X2_26/A OAI21X1_599/B gnd INVX1_232/A vdd AOI21X1
XAOI21X1_206 BUFX4_114/Y OAI22X1_32/D OAI21X1_550/Y gnd OAI21X1_551/C vdd AOI21X1
XAOI21X1_228 NAND2X1_498/Y AOI21X1_228/B OAI22X1_35/A gnd OAI21X1_581/A vdd AOI21X1
XAOI22X1_22 BUFX4_56/Y INVX1_219/A BUFX4_4/Y INVX1_223/Y gnd AOI22X1_22/Y vdd AOI22X1
XAOI22X1_11 BUFX4_153/Y NOR2X1_202/B BUFX4_58/Y INVX1_169/A gnd AOI22X1_11/Y vdd AOI22X1
XAOI22X1_55 INVX8_17/A NOR2X1_41/Y NAND2X1_52/Y BUFX4_3/Y gnd AOI22X1_55/Y vdd AOI22X1
XAOI22X1_33 BUFX4_150/Y NOR2X1_17/Y XOR2X1_7/Y INVX8_14/A gnd NAND3X1_57/C vdd AOI22X1
XAOI22X1_44 BUFX4_60/Y NAND3X1_1/A NAND2X1_43/Y BUFX4_1/Y gnd AOI22X1_44/Y vdd AOI22X1
XFILL_23_1_0 gnd vdd FILL
XOAI22X1_6 BUFX4_86/Y OAI22X1_6/B OAI22X1_6/C OR2X2_40/B gnd OAI22X1_6/Y vdd OAI22X1
XFILL_6_2_0 gnd vdd FILL
XFILL_14_1_0 gnd vdd FILL
XFILL_33_1 gnd vdd FILL
XNOR2X1_412 INVX1_199/A NOR2X1_412/B gnd NOR2X1_412/Y vdd NOR2X1
XNOR2X1_423 NOR2X1_423/A NOR2X1_423/B gnd NOR2X1_423/Y vdd NOR2X1
XNOR2X1_467 BUFX4_83/Y NOR2X1_467/B gnd NOR2X1_467/Y vdd NOR2X1
XNOR2X1_401 OR2X2_48/B BUFX2_23/A gnd NOR2X1_401/Y vdd NOR2X1
XNOR2X1_456 BUFX4_114/Y NOR2X1_456/B gnd NOR2X1_456/Y vdd NOR2X1
XNOR2X1_434 BUFX4_97/Y BUFX2_6/A gnd NOR2X1_434/Y vdd NOR2X1
XNOR2X1_445 BUFX4_100/Y BUFX2_9/A gnd NOR2X1_445/Y vdd NOR2X1
XOAI21X1_929 BUFX4_158/Y XNOR2X1_27/Y BUFX4_99/Y gnd NOR2X1_500/A vdd OAI21X1
XOAI21X1_918 BUFX4_96/Y XNOR2X1_47/Y OAI21X1_918/C gnd OAI21X1_919/A vdd OAI21X1
XOAI21X1_907 XNOR2X1_46/B OAI21X1_907/B OAI21X1_907/C gnd AOI22X1_54/D vdd OAI21X1
XNOR2X1_478 BUFX4_83/Y NOR2X1_478/B gnd NOR2X1_478/Y vdd NOR2X1
XNOR2X1_489 NOR2X1_489/A NOR2X1_489/B gnd NOR2X1_489/Y vdd NOR2X1
XINVX2_15 operand_A[15] gnd INVX2_15/Y vdd INVX2
XINVX2_26 operand_A[8] gnd INVX2_26/Y vdd INVX2
XINVX2_59 INVX2_59/A gnd OR2X2_9/B vdd INVX2
XINVX2_37 alu_op[1] gnd INVX2_37/Y vdd INVX2
XINVX2_48 INVX2_48/A gnd INVX2_48/Y vdd INVX2
XFILL_30_4_1 gnd vdd FILL
XNAND2X1_209 MUX2X1_98/S INVX1_48/Y gnd OAI21X1_176/C vdd NAND2X1
XNOR2X1_286 AND2X2_32/Y NOR2X1_286/B gnd NOR2X1_286/Y vdd NOR2X1
XNOR2X1_275 BUFX4_102/Y BUFX2_54/A gnd NOR2X1_275/Y vdd NOR2X1
XNOR2X1_242 INVX2_42/Y INVX1_197/Y gnd INVX1_201/A vdd NOR2X1
XNOR2X1_297 INVX1_229/A AND2X2_35/Y gnd INVX2_79/A vdd NOR2X1
XNOR2X1_264 OR2X2_30/B OR2X2_30/A gnd NOR2X1_264/Y vdd NOR2X1
XNOR2X1_220 INVX2_75/Y NOR2X1_220/B gnd NOR2X1_226/B vdd NOR2X1
XNOR2X1_231 NOR2X1_231/A NOR2X1_231/B gnd INVX1_186/A vdd NOR2X1
XBUFX4_171 INVX8_10/Y gnd BUFX4_171/Y vdd BUFX4
XNOR2X1_253 NOR2X1_253/A OAI22X1_28/A gnd NOR2X1_253/Y vdd NOR2X1
XBUFX4_193 operand_B[1] gnd MUX2X1_97/S vdd BUFX4
XBUFX4_182 operand_B[4] gnd NOR2X1_75/A vdd BUFX4
XBUFX4_160 INVX8_5/Y gnd MUX2X1_32/S vdd BUFX4
XFILL_21_4_1 gnd vdd FILL
XOAI21X1_704 INVX4_8/Y MUX2X1_6/S OAI21X1_704/C gnd OAI21X1_704/Y vdd OAI21X1
XOAI21X1_726 INVX1_293/Y MUX2X1_71/S OAI21X1_726/C gnd MUX2X1_120/A vdd OAI21X1
XOAI21X1_715 NOR2X1_431/Y AOI21X1_75/B BUFX4_111/Y gnd OAI21X1_715/Y vdd OAI21X1
XOAI21X1_759 XNOR2X1_20/Y OAI21X1_759/B OAI21X1_759/C gnd NAND3X1_61/A vdd OAI21X1
XOAI21X1_737 INVX1_295/Y BUFX4_125/Y OAI21X1_737/C gnd OAI21X1_738/B vdd OAI21X1
XOAI21X1_748 BUFX4_24/Y NOR2X1_464/B OAI21X1_748/C gnd MUX2X1_107/A vdd OAI21X1
XFILL_29_5_1 gnd vdd FILL
XFILL_28_0_0 gnd vdd FILL
XFILL_3_0_0 gnd vdd FILL
XFILL_4_5_1 gnd vdd FILL
XFILL_12_4_1 gnd vdd FILL
XINVX8_2 INVX8_2/A gnd INVX8_2/Y vdd INVX8
XBUFX4_44 operand_B[0] gnd MUX2X1_4/S vdd BUFX4
XBUFX4_55 operand_B[0] gnd MUX2X1_8/S vdd BUFX4
XBUFX4_66 INVX8_1/Y gnd BUFX4_66/Y vdd BUFX4
XBUFX4_33 operand_B[3] gnd INVX8_2/A vdd BUFX4
XBUFX4_11 INVX8_19/Y gnd BUFX4_11/Y vdd BUFX4
XBUFX4_77 INVX8_4/Y gnd BUFX4_77/Y vdd BUFX4
XBUFX4_22 INVX8_2/Y gnd BUFX4_22/Y vdd BUFX4
XBUFX4_99 DFFSR_1/Q gnd BUFX4_99/Y vdd BUFX4
XFILL_19_0_0 gnd vdd FILL
XBUFX4_88 BUFX4_91/A gnd INVX8_12/A vdd BUFX4
XOR2X2_14 OR2X2_14/A OR2X2_19/B gnd OR2X2_14/Y vdd OR2X2
XOR2X2_36 OR2X2_36/A OR2X2_36/B gnd OR2X2_36/Y vdd OR2X2
XOR2X2_25 OR2X2_25/A OR2X2_25/B gnd OR2X2_25/Y vdd OR2X2
XOR2X2_47 OR2X2_47/A OR2X2_47/B gnd OR2X2_47/Y vdd OR2X2
XXNOR2X1_9 operand_A[8] operand_B[8] gnd INVX1_17/A vdd XNOR2X1
XOR2X2_7 OR2X2_7/A OR2X2_7/B gnd OR2X2_7/Y vdd OR2X2
XOAI21X1_501 INVX1_204/A OAI21X1_501/B OAI21X1_501/C gnd OAI21X1_501/Y vdd OAI21X1
XOAI21X1_512 INVX1_205/Y BUFX4_70/Y OAI21X1_512/C gnd OAI21X1_558/B vdd OAI21X1
XINVX1_9 operand_B[22] gnd INVX1_9/Y vdd INVX1
XOAI21X1_523 AOI21X1_86/Y BUFX4_179/Y INVX4_11/Y gnd OAI21X1_523/Y vdd OAI21X1
XINVX8_14 INVX8_14/A gnd INVX8_14/Y vdd INVX8
XOAI21X1_545 INVX1_222/A INVX1_223/A NOR2X1_293/Y gnd OAI21X1_546/C vdd OAI21X1
XOAI21X1_589 AND2X2_41/Y NOR2X1_341/A INVX2_86/Y gnd NAND3X1_35/B vdd OAI21X1
XOAI21X1_556 INVX2_80/Y BUFX4_46/Y OAI21X1_556/C gnd OAI21X1_577/B vdd OAI21X1
XOAI21X1_534 INVX2_53/Y MUX2X1_4/S OAI21X1_534/C gnd INVX1_220/A vdd OAI21X1
XOAI21X1_567 INVX2_39/Y MUX2X1_5/S OAI21X1_63/C gnd MUX2X1_56/B vdd OAI21X1
XOAI21X1_578 MUX2X1_62/B BUFX4_136/Y OAI21X1_578/C gnd MUX2X1_55/B vdd OAI21X1
XNAND2X1_540 operand_B[28] INVX4_2/Y gnd NOR2X1_414/A vdd NAND2X1
XNAND2X1_551 operand_B[45] INVX4_14/Y gnd OAI21X1_669/C vdd NAND2X1
XNAND2X1_584 BUFX4_72/Y OAI21X1_676/Y gnd OAI21X1_725/C vdd NAND2X1
XNAND2X1_562 MUX2X1_8/S operand_A[13] gnd OAI21X1_685/C vdd NAND2X1
XNAND2X1_595 BUFX4_133/Y INVX1_287/A gnd OAI21X1_747/C vdd NAND2X1
XNAND2X1_573 BUFX4_133/Y OAI21X1_708/Y gnd OAI21X1_711/C vdd NAND2X1
XFILL_9_2 gnd vdd FILL
XFILL_26_3_1 gnd vdd FILL
XFILL_1_3_1 gnd vdd FILL
XOAI21X1_331 INVX1_144/Y NOR2X1_420/A NOR2X1_183/A gnd OR2X2_12/A vdd OAI21X1
XOAI21X1_364 BUFX4_61/Y INVX1_156/Y OAI21X1_364/C gnd OAI21X1_364/Y vdd OAI21X1
XOAI21X1_342 BUFX4_21/Y INVX1_55/Y OR2X2_13/Y gnd OAI21X1_342/Y vdd OAI21X1
XOAI21X1_320 INVX1_137/Y BUFX4_39/Y OAI21X1_320/C gnd INVX1_138/A vdd OAI21X1
XOAI21X1_353 INVX1_150/Y MUX2X1_49/S OAI21X1_353/C gnd OAI21X1_353/Y vdd OAI21X1
XAND2X2_9 AND2X2_9/A NOR2X1_3/Y gnd AND2X2_9/Y vdd AND2X2
XOAI21X1_386 NOR2X1_194/Y NOR2X1_193/Y BUFX4_84/Y gnd NAND3X1_18/A vdd OAI21X1
XOAI21X1_397 OAI21X1_397/A INVX8_2/A OAI21X1_397/C gnd OAI22X1_16/A vdd OAI21X1
XOAI21X1_375 BUFX4_23/Y OAI21X1_375/B OAI21X1_375/C gnd OAI21X1_375/Y vdd OAI21X1
XFILL_9_4_1 gnd vdd FILL
XNAND2X1_392 BUFX4_134/Y OAI21X1_349/Y gnd OAI21X1_414/C vdd NAND2X1
XNAND2X1_370 MUX2X1_62/S OAI21X1_372/Y gnd OAI21X1_373/C vdd NAND2X1
XNAND2X1_381 BUFX4_22/Y OAI21X1_228/A gnd OAI21X1_390/C vdd NAND2X1
XFILL_17_3_1 gnd vdd FILL
XINVX1_225 INVX1_225/A gnd INVX1_225/Y vdd INVX1
XINVX1_203 operand_B[49] gnd INVX1_203/Y vdd INVX1
XINVX1_214 INVX1_214/A gnd INVX1_214/Y vdd INVX1
XOAI21X1_172 INVX2_1/Y operand_A[29] AND2X2_2/A gnd OAI21X1_173/A vdd OAI21X1
XOAI21X1_150 OAI21X1_150/A INVX1_2/A AOI21X1_45/Y gnd AOI21X1_46/C vdd OAI21X1
XAOI22X1_4 BUFX4_148/Y INVX4_15/Y AOI22X1_4/C BUFX4_57/Y gnd AOI22X1_4/Y vdd AOI22X1
XOAI21X1_183 XOR2X1_3/A OAI21X1_82/Y OAI21X1_183/C gnd OAI21X1_183/Y vdd OAI21X1
XOAI21X1_161 NOR2X1_117/Y OAI21X1_806/C OAI21X1_639/C gnd AOI21X1_53/A vdd OAI21X1
XOAI21X1_194 INVX1_91/Y BUFX4_67/Y OAI21X1_194/C gnd INVX1_92/A vdd OAI21X1
XINVX1_247 INVX1_247/A gnd INVX1_247/Y vdd INVX1
XINVX1_236 INVX1_236/A gnd INVX1_236/Y vdd INVX1
XINVX1_258 INVX1_258/A gnd INVX1_258/Y vdd INVX1
XINVX1_269 BUFX2_3/A gnd INVX1_269/Y vdd INVX1
XNAND2X1_14 operand_B[21] operand_A[21] gnd OAI21X1_4/C vdd NAND2X1
XNAND2X1_25 OR2X2_43/B INVX4_7/Y gnd INVX2_92/A vdd NAND2X1
XNAND2X1_47 AOI22X1_1/A NAND2X1_47/B gnd NOR2X1_67/A vdd NAND2X1
XNAND2X1_58 NAND2X1_58/A NAND2X1_58/B gnd NAND2X1_59/B vdd NAND2X1
XNAND2X1_36 NAND2X1_36/A NAND2X1_36/B gnd XNOR2X1_41/B vdd NAND2X1
XNAND2X1_69 XNOR2X1_16/Y XNOR2X1_17/Y gnd OAI21X1_28/A vdd NAND2X1
XFILL_32_1_1 gnd vdd FILL
XAOI21X1_207 NAND2X1_476/Y AOI21X1_207/B OAI21X1_551/Y gnd AOI21X1_208/B vdd AOI21X1
XAOI22X1_23 BUFX4_56/Y INVX2_79/A BUFX4_4/Y INVX1_229/Y gnd NAND3X1_33/B vdd AOI22X1
XAOI21X1_218 OAI21X1_660/C INVX1_226/A NOR2X1_313/Y gnd NAND2X1_492/A vdd AOI21X1
XAOI21X1_229 NOR2X1_22/A OAI22X1_35/D OAI21X1_580/Y gnd OAI21X1_581/C vdd AOI21X1
XAOI22X1_12 AOI22X1_12/A INVX4_20/A INVX8_18/A AND2X2_59/A gnd NAND3X1_20/C vdd AOI22X1
XAOI22X1_56 BUFX4_13/Y INVX1_275/Y NOR2X1_501/Y AOI22X1_56/D gnd AOI22X1_56/Y vdd
+ AOI22X1
XAOI22X1_34 BUFX4_14/Y INVX1_267/Y OAI22X1_27/Y NOR2X1_441/Y gnd DFFPOSX1_5/D vdd
+ AOI22X1
XAOI22X1_45 BUFX4_15/Y INVX1_273/Y AND2X2_68/Y AND2X2_67/Y gnd AOI22X1_45/Y vdd AOI22X1
XFILL_23_1_1 gnd vdd FILL
XOAI22X1_7 OAI22X1_9/A OR2X2_21/B OAI22X1_7/C OAI22X1_7/D gnd OAI22X1_7/Y vdd OAI22X1
XFILL_6_2_1 gnd vdd FILL
XFILL_14_1_1 gnd vdd FILL
XFILL_33_2 gnd vdd FILL
XFILL_26_1 gnd vdd FILL
XNOR2X1_424 NOR2X1_424/A NOR2X1_424/B gnd NOR2X1_424/Y vdd NOR2X1
XNOR2X1_413 NOR2X1_413/A NOR2X1_413/B gnd NOR2X1_413/Y vdd NOR2X1
XNOR2X1_435 BUFX4_172/Y NOR2X1_435/B gnd NOR2X1_435/Y vdd NOR2X1
XNOR2X1_457 INVX1_17/A AOI21X1_9/Y gnd INVX1_306/A vdd NOR2X1
XNOR2X1_479 NOR2X1_479/A NOR2X1_479/B gnd NOR2X1_479/Y vdd NOR2X1
XNOR2X1_402 BUFX2_18/A BUFX2_17/A gnd NOR2X1_402/Y vdd NOR2X1
XNOR2X1_446 MUX2X1_32/S NOR2X1_446/B gnd NOR2X1_447/B vdd NOR2X1
XNOR2X1_468 NOR2X1_468/A NOR2X1_468/B gnd NOR2X1_468/Y vdd NOR2X1
XOAI21X1_919 OAI21X1_919/A OAI21X1_919/B BUFX4_99/Y gnd OAI21X1_920/C vdd OAI21X1
XOAI21X1_908 MUX2X1_57/S NOR2X1_449/B OAI21X1_908/C gnd OAI21X1_908/Y vdd OAI21X1
XINVX2_38 operand_A[54] gnd INVX2_38/Y vdd INVX2
XINVX2_49 INVX2_49/A gnd INVX2_49/Y vdd INVX2
XINVX2_27 operand_A[11] gnd INVX2_27/Y vdd INVX2
XINVX2_16 operand_A[14] gnd INVX2_16/Y vdd INVX2
XCLKBUF1_1 clk gnd CLKBUF1_1/Y vdd CLKBUF1
XBUFX4_172 INVX8_10/Y gnd BUFX4_172/Y vdd BUFX4
XBUFX4_161 INVX8_5/Y gnd NOR2X1_80/A vdd BUFX4
XBUFX4_150 NOR2X1_89/Y gnd BUFX4_150/Y vdd BUFX4
XNOR2X1_276 operand_A[52] operand_B[52] gnd OAI22X1_11/D vdd NOR2X1
XNOR2X1_243 INVX1_202/A INVX1_201/A gnd AND2X2_26/B vdd NOR2X1
XNOR2X1_265 AND2X2_26/B INVX1_204/A gnd NOR2X1_265/Y vdd NOR2X1
XNOR2X1_298 operand_B[54] INVX2_38/Y gnd INVX1_226/A vdd NOR2X1
XNOR2X1_210 OAI22X1_7/D NOR2X1_210/B gnd INVX2_74/A vdd NOR2X1
XNOR2X1_221 BUFX4_27/Y NOR2X1_226/B gnd NOR2X1_221/Y vdd NOR2X1
XNOR2X1_232 operand_B[44] INVX2_46/Y gnd NOR2X1_232/Y vdd NOR2X1
XNOR2X1_254 OR2X2_8/B NOR2X1_254/B gnd NOR2X1_254/Y vdd NOR2X1
XOAI21X1_705 BUFX4_72/Y MUX2X1_78/Y OAI21X1_705/C gnd OAI21X1_762/B vdd OAI21X1
XNOR2X1_287 INVX8_7/Y MUX2X1_49/Y gnd NOR2X1_287/Y vdd NOR2X1
XBUFX4_194 operand_B[1] gnd MUX2X1_98/S vdd BUFX4
XBUFX4_183 operand_B[4] gnd BUFX4_183/Y vdd BUFX4
XOAI21X1_749 INVX1_296/Y BUFX4_171/Y BUFX4_113/Y gnd OAI22X1_27/C vdd OAI21X1
XOAI21X1_716 INVX1_285/Y BUFX4_76/Y OAI21X1_716/C gnd INVX1_291/A vdd OAI21X1
XOAI21X1_738 INVX8_2/A OAI21X1_738/B OR2X2_39/Y gnd INVX1_318/A vdd OAI21X1
XOAI21X1_727 OAI21X1_727/A BUFX4_42/Y OAI21X1_727/C gnd MUX2X1_124/A vdd OAI21X1
XFILL_28_0_1 gnd vdd FILL
XFILL_3_0_1 gnd vdd FILL
XINVX8_3 INVX8_3/A gnd INVX8_3/Y vdd INVX8
XAOI21X1_390 XNOR2X1_46/B OAI21X1_907/B BUFX4_96/Y gnd OAI21X1_907/C vdd AOI21X1
XBUFX4_56 BUFX4_60/A gnd BUFX4_56/Y vdd BUFX4
XFILL_19_0_1 gnd vdd FILL
XBUFX4_12 INVX8_19/Y gnd BUFX4_12/Y vdd BUFX4
XBUFX4_45 operand_B[0] gnd MUX2X1_9/S vdd BUFX4
XBUFX4_34 operand_B[3] gnd XOR2X1_4/A vdd BUFX4
XBUFX4_67 INVX8_1/Y gnd BUFX4_67/Y vdd BUFX4
XBUFX4_23 INVX8_2/Y gnd BUFX4_23/Y vdd BUFX4
XBUFX4_78 INVX8_4/Y gnd BUFX4_78/Y vdd BUFX4
XBUFX4_89 BUFX4_91/A gnd BUFX4_89/Y vdd BUFX4
XOR2X2_37 OR2X2_37/A OR2X2_37/B gnd OR2X2_37/Y vdd OR2X2
XOR2X2_26 OR2X2_26/A OR2X2_8/B gnd OR2X2_26/Y vdd OR2X2
XOR2X2_15 OR2X2_15/A OR2X2_19/B gnd OR2X2_15/Y vdd OR2X2
XOR2X2_48 OR2X2_48/A OR2X2_48/B gnd OR2X2_48/Y vdd OR2X2
XOR2X2_8 OR2X2_8/A OR2X2_8/B gnd OR2X2_8/Y vdd OR2X2
XOAI21X1_546 INVX2_53/Y operand_B[53] OAI21X1_546/C gnd OAI21X1_546/Y vdd OAI21X1
XOAI21X1_535 INVX1_220/Y MUX2X1_23/S OAI21X1_535/C gnd OAI21X1_535/Y vdd OAI21X1
XOAI21X1_557 INVX1_220/Y BUFX4_70/Y OAI21X1_557/C gnd INVX1_227/A vdd OAI21X1
XOAI21X1_513 INVX1_213/Y MUX2X1_66/S OAI21X1_513/C gnd MUX2X1_58/B vdd OAI21X1
XOAI21X1_524 BUFX4_163/Y INVX1_132/Y OAI21X1_524/C gnd MUX2X1_48/B vdd OAI21X1
XOAI21X1_502 INVX1_209/Y MUX2X1_64/S INVX8_7/A gnd OAI21X1_502/Y vdd OAI21X1
XINVX8_15 INVX8_15/A gnd INVX8_15/Y vdd INVX8
XOAI21X1_579 operand_A[57] operand_B[57] BUFX4_4/Y gnd AND2X2_39/B vdd OAI21X1
XOAI21X1_568 BUFX4_134/Y MUX2X1_60/B OAI21X1_568/C gnd MUX2X1_54/B vdd OAI21X1
XNAND2X1_530 NOR2X1_378/Y NOR2X1_379/Y gnd NOR2X1_380/B vdd NAND2X1
XNAND2X1_541 operand_B[49] INVX2_52/Y gnd OAI21X1_659/C vdd NAND2X1
XNAND2X1_552 operand_B[44] INVX2_46/Y gnd OAI21X1_669/B vdd NAND2X1
XNAND2X1_585 MUX2X1_71/S MUX2X1_111/B gnd OAI21X1_726/C vdd NAND2X1
XNAND2X1_563 XOR2X1_3/A OAI21X1_686/Y gnd OAI21X1_687/C vdd NAND2X1
XNAND2X1_574 MUX2X1_97/S MUX2X1_80/Y gnd OAI21X1_710/C vdd NAND2X1
XNAND2X1_596 BUFX4_24/Y OAI21X1_747/Y gnd OAI21X1_748/C vdd NAND2X1
XOAI21X1_354 OAI22X1_9/A INVX1_148/A OAI21X1_354/C gnd NOR2X1_175/B vdd OAI21X1
XOAI21X1_332 INVX1_146/Y BUFX4_16/Y OAI21X1_332/C gnd AND2X2_14/A vdd OAI21X1
XOAI21X1_398 OAI22X1_16/A INVX8_8/Y INVX8_15/Y gnd OAI21X1_404/C vdd OAI21X1
XOAI21X1_365 BUFX4_25/Y OAI21X1_365/B OAI21X1_365/C gnd MUX2X1_126/A vdd OAI21X1
XOAI21X1_376 NOR2X1_316/B OR2X2_43/B OAI21X1_376/C gnd OAI21X1_377/A vdd OAI21X1
XOAI21X1_387 INVX1_166/Y MUX2X1_99/S BUFX4_38/Y gnd OAI21X1_388/C vdd OAI21X1
XOAI21X1_321 INVX1_104/Y MUX2X1_27/S OAI21X1_321/C gnd INVX1_139/A vdd OAI21X1
XOAI21X1_343 BUFX4_173/Y OAI21X1_780/A OAI22X1_6/Y gnd NOR2X1_171/B vdd OAI21X1
XOAI21X1_310 BUFX4_22/Y INVX1_183/A OAI21X1_310/C gnd MUX2X1_34/B vdd OAI21X1
XNAND2X1_382 INVX1_154/A INVX1_162/A gnd NOR2X1_219/A vdd NAND2X1
XNAND2X1_371 BUFX4_18/Y INVX1_160/Y gnd OAI21X1_374/C vdd NAND2X1
XNAND2X1_393 BUFX4_25/Y INVX1_175/Y gnd OAI21X1_415/C vdd NAND2X1
XNAND2X1_360 MUX2X1_49/S NOR2X1_300/B gnd OAI21X1_353/C vdd NAND2X1
XINVX1_215 BUFX2_55/A gnd INVX1_215/Y vdd INVX1
XINVX1_204 INVX1_204/A gnd INVX1_204/Y vdd INVX1
XINVX1_226 INVX1_226/A gnd INVX1_226/Y vdd INVX1
XOAI21X1_173 OAI21X1_173/A NOR2X1_121/B AOI21X1_59/Y gnd AOI21X1_60/C vdd OAI21X1
XINVX1_248 INVX1_248/A gnd INVX1_248/Y vdd INVX1
XINVX1_237 INVX1_237/A gnd INVX1_237/Y vdd INVX1
XINVX1_259 INVX1_259/A gnd INVX1_259/Y vdd INVX1
XOAI21X1_151 INVX1_10/A NOR2X1_106/B AOI21X1_46/Y gnd AOI21X1_47/C vdd OAI21X1
XOAI21X1_140 INVX2_55/Y BUFX4_46/Y OAI21X1_348/C gnd OAI21X1_140/Y vdd OAI21X1
XAOI22X1_5 BUFX4_57/Y INVX4_16/Y BUFX4_3/Y OR2X2_6/Y gnd AOI22X1_5/Y vdd AOI22X1
XOAI21X1_184 MUX2X1_30/S OAI21X1_299/B OAI21X1_184/C gnd INVX1_88/A vdd OAI21X1
XOAI21X1_162 NOR2X1_118/Y OAI21X1_162/B INVX1_83/Y gnd AOI21X1_53/C vdd OAI21X1
XOAI21X1_195 INVX1_93/Y BUFX4_67/Y OAI21X1_195/C gnd INVX1_128/A vdd OAI21X1
XFILL_10_5_0 gnd vdd FILL
XNAND2X1_48 operand_A[26] INVX1_22/Y gnd OAI21X1_33/C vdd NAND2X1
XNAND2X1_59 NAND2X1_59/A NAND2X1_59/B gnd OR2X2_2/B vdd NAND2X1
XNAND2X1_15 INVX2_8/Y INVX1_8/Y gnd AOI21X1_4/A vdd NAND2X1
XNAND2X1_37 operand_A[12] INVX1_19/Y gnd NAND2X1_39/A vdd NAND2X1
XNAND2X1_26 NAND2X1_26/A INVX2_92/A gnd NAND3X1_4/B vdd NAND2X1
XNAND2X1_190 operand_A[32] operand_B[32] gnd INVX4_15/A vdd NAND2X1
XAOI21X1_208 OAI21X1_544/Y AOI21X1_208/B NOR2X1_295/Y gnd DFFPOSX1_55/D vdd AOI21X1
XAOI21X1_219 INVX2_81/Y OAI21X1_566/B BUFX4_94/Y gnd OAI21X1_566/C vdd AOI21X1
XAOI22X1_24 BUFX4_149/Y NOR2X1_321/A BUFX4_56/Y INVX2_81/A gnd AND2X2_37/A vdd AOI22X1
XAOI22X1_57 BUFX4_13/Y INVX1_274/Y AOI22X1_57/C AOI22X1_57/D gnd AOI22X1_57/Y vdd
+ AOI22X1
XAOI22X1_13 INVX8_17/A AND2X2_21/Y BUFX4_57/Y INVX2_75/A gnd AOI22X1_13/Y vdd AOI22X1
XAOI22X1_35 INVX8_14/A NAND3X1_4/A INVX1_301/Y BUFX4_2/Y gnd NAND3X1_62/B vdd AOI22X1
XAOI22X1_46 BUFX4_152/Y NOR2X1_7/Y AOI21X1_2/A BUFX4_3/Y gnd AND2X2_70/A vdd AOI22X1
XOAI22X1_8 OR2X2_19/B OAI22X1_8/B OAI22X1_8/C OAI22X1_8/D gnd OR2X2_27/B vdd OAI22X1
XAOI21X1_90 INVX2_65/A AOI21X1_90/B BUFX4_28/Y gnd AOI21X1_90/Y vdd AOI21X1
XFILL_26_2 gnd vdd FILL
XNOR2X1_414 NOR2X1_414/A NAND2X1_3/Y gnd NOR2X1_414/Y vdd NOR2X1
XFILL_19_1 gnd vdd FILL
XNOR2X1_403 NOR2X1_403/A NOR2X1_403/B gnd NOR2X1_403/Y vdd NOR2X1
XNOR2X1_425 NOR2X1_19/B MUX2X1_76/Y gnd NOR2X1_425/Y vdd NOR2X1
XNOR2X1_436 INVX8_15/Y OR2X2_10/Y gnd NOR2X1_437/B vdd NOR2X1
XNOR2X1_469 BUFX4_100/Y BUFX2_16/A gnd NOR2X1_469/Y vdd NOR2X1
XNOR2X1_458 MUX2X1_25/S NOR2X1_458/B gnd NOR2X1_458/Y vdd NOR2X1
XNOR2X1_447 INVX8_4/A NOR2X1_447/B gnd NOR2X1_447/Y vdd NOR2X1
XOAI21X1_909 OAI21X1_23/A XNOR2X1_29/Y OAI21X1_909/C gnd OAI21X1_909/Y vdd OAI21X1
XINVX2_39 operand_A[56] gnd INVX2_39/Y vdd INVX2
XINVX2_17 INVX2_17/A gnd INVX2_17/Y vdd INVX2
XINVX2_28 operand_B[11] gnd INVX2_28/Y vdd INVX2
XFILL_24_4_0 gnd vdd FILL
XFILL_7_5_0 gnd vdd FILL
XFILL_15_4_0 gnd vdd FILL
XMUX2X1_1 operand_A[1] operand_A[2] MUX2X1_1/S gnd MUX2X1_1/Y vdd MUX2X1
XCLKBUF1_2 clk gnd CLKBUF1_2/Y vdd CLKBUF1
XNOR2X1_200 INVX2_71/Y INVX2_72/Y gnd NOR2X1_202/B vdd NOR2X1
XBUFX4_151 NOR2X1_89/Y gnd INVX8_17/A vdd BUFX4
XNOR2X1_233 operand_B[45] INVX4_14/Y gnd NOR2X1_233/Y vdd NOR2X1
XNOR2X1_222 BUFX4_41/Y NOR2X1_222/B gnd INVX1_176/A vdd NOR2X1
XBUFX4_140 NOR2X1_72/Y gnd BUFX4_140/Y vdd BUFX4
XBUFX4_173 INVX8_18/Y gnd BUFX4_173/Y vdd BUFX4
XBUFX4_195 operand_B[1] gnd NOR2X1_82/A vdd BUFX4
XBUFX4_184 operand_B[4] gnd BUFX4_184/Y vdd BUFX4
XBUFX4_162 INVX8_5/Y gnd BUFX4_162/Y vdd BUFX4
XNOR2X1_211 MUX2X1_32/S OAI22X1_19/C gnd NOR2X1_211/Y vdd NOR2X1
XNOR2X1_255 BUFX4_102/Y BUFX2_52/A gnd NOR2X1_255/Y vdd NOR2X1
XNOR2X1_277 OAI22X1_11/D AND2X2_32/Y gnd INVX2_78/A vdd NOR2X1
XNOR2X1_244 NOR2X1_244/A OR2X2_28/A gnd NOR2X1_244/Y vdd NOR2X1
XNOR2X1_288 OR2X2_8/B NOR2X1_288/B gnd NOR2X1_288/Y vdd NOR2X1
XNOR2X1_266 BUFX4_25/Y MUX2X1_38/B gnd NOR2X1_266/Y vdd NOR2X1
XNOR2X1_299 BUFX4_79/Y NOR2X1_497/B gnd NOR2X1_299/Y vdd NOR2X1
XOAI21X1_717 INVX1_288/Y BUFX4_74/Y OAI21X1_717/C gnd MUX2X1_110/B vdd OAI21X1
XOAI21X1_739 MUX2X1_23/S MUX2X1_90/B OAI21X1_739/C gnd MUX2X1_114/B vdd OAI21X1
XOAI21X1_728 MUX2X1_124/A BUFX4_162/Y AND2X2_11/B gnd OAI21X1_728/Y vdd OAI21X1
XOAI21X1_706 MUX2X1_51/S OAI21X1_762/B OAI21X1_706/C gnd MUX2X1_118/A vdd OAI21X1
XAOI21X1_380 NOR2X1_66/Y OAI21X1_32/Y OAI21X1_26/Y gnd OAI21X1_901/A vdd AOI21X1
XAOI21X1_391 BUFX4_79/Y OAI21X1_908/Y INVX8_9/Y gnd OAI22X1_33/C vdd AOI21X1
XINVX8_4 INVX8_4/A gnd INVX8_4/Y vdd INVX8
XBUFX4_57 BUFX4_60/A gnd BUFX4_57/Y vdd BUFX4
XBUFX4_68 INVX8_1/Y gnd BUFX4_68/Y vdd BUFX4
XBUFX4_13 INVX8_19/Y gnd BUFX4_13/Y vdd BUFX4
XBUFX4_79 INVX8_4/Y gnd BUFX4_79/Y vdd BUFX4
XBUFX4_46 operand_B[0] gnd BUFX4_46/Y vdd BUFX4
XBUFX4_35 operand_B[3] gnd BUFX4_35/Y vdd BUFX4
XBUFX4_24 INVX8_2/Y gnd BUFX4_24/Y vdd BUFX4
XFILL_30_2_0 gnd vdd FILL
XOR2X2_9 OR2X2_9/A OR2X2_9/B gnd OR2X2_9/Y vdd OR2X2
XOR2X2_38 OR2X2_38/A OR2X2_38/B gnd OR2X2_38/Y vdd OR2X2
XOR2X2_49 OR2X2_49/A OR2X2_49/B gnd OR2X2_49/Y vdd OR2X2
XOR2X2_27 OR2X2_27/A OR2X2_27/B gnd OR2X2_27/Y vdd OR2X2
XOR2X2_16 OR2X2_16/A OR2X2_16/B gnd OR2X2_16/Y vdd OR2X2
XINVX8_16 BUFX4_5/Y gnd INVX8_16/Y vdd INVX8
XOAI21X1_503 INVX2_41/Y BUFX4_53/Y OAI21X1_70/C gnd INVX1_210/A vdd OAI21X1
XOAI21X1_525 INVX2_40/Y MUX2X1_8/S OAI21X1_68/C gnd MUX2X1_50/B vdd OAI21X1
XOAI21X1_547 INVX2_38/Y MUX2X1_9/S OAI21X1_67/C gnd MUX2X1_53/B vdd OAI21X1
XFILL_21_2_0 gnd vdd FILL
XOAI21X1_569 NOR2X1_316/Y NOR2X1_315/Y INVX8_7/A gnd OAI21X1_569/Y vdd OAI21X1
XOAI21X1_536 INVX1_206/Y MUX2X1_66/S OAI21X1_536/C gnd MUX2X1_63/A vdd OAI21X1
XOAI21X1_558 MUX2X1_62/S OAI21X1_558/B OAI21X1_558/C gnd OAI21X1_631/A vdd OAI21X1
XOAI21X1_514 INVX1_175/Y BUFX4_17/Y OAI21X1_514/C gnd MUX2X1_46/A vdd OAI21X1
XNAND2X1_520 NOR2X1_80/A NOR2X1_228/Y gnd OAI21X1_946/A vdd NAND2X1
XNAND2X1_531 NOR2X1_382/Y NOR2X1_383/Y gnd NOR2X1_384/B vdd NAND2X1
XFILL_29_3_0 gnd vdd FILL
XNAND2X1_542 operand_B[48] INVX2_42/Y gnd OAI21X1_659/B vdd NAND2X1
XNAND2X1_553 operand_B[41] INVX2_54/Y gnd OAI21X1_672/C vdd NAND2X1
XNAND2X1_564 NOR2X1_83/A MUX2X1_106/A gnd OAI21X1_688/C vdd NAND2X1
XFILL_4_3_0 gnd vdd FILL
XNAND2X1_597 OAI21X1_752/Y NOR2X1_440/Y gnd NOR2X1_441/B vdd NAND2X1
XNAND2X1_575 OR2X2_39/B MUX2X1_119/A gnd NAND2X1_575/Y vdd NAND2X1
XNAND2X1_586 BUFX4_41/Y MUX2X1_120/A gnd OAI21X1_727/C vdd NAND2X1
XFILL_12_2_0 gnd vdd FILL
XOAI21X1_344 OAI21X1_344/A NAND3X1_13/Y BUFX4_101/Y gnd OAI21X1_345/C vdd OAI21X1
XOAI21X1_322 INVX2_55/Y BUFX4_48/Y OAI21X1_322/C gnd INVX1_140/A vdd OAI21X1
XOAI21X1_300 BUFX4_133/Y MUX2X1_24/B OAI21X1_300/C gnd MUX2X1_33/B vdd OAI21X1
XOAI21X1_333 BUFX4_21/Y INVX1_53/Y OR2X2_13/Y gnd OAI21X1_333/Y vdd OAI21X1
XOAI21X1_366 NOR2X1_80/A NOR2X1_317/B OAI21X1_366/C gnd AND2X2_57/A vdd OAI21X1
XOAI21X1_355 NAND3X1_14/Y OR2X2_32/B NOR2X1_175/Y gnd OAI21X1_355/Y vdd OAI21X1
XOAI21X1_377 OAI21X1_377/A BUFX4_116/Y OAI21X1_377/C gnd NAND3X1_17/B vdd OAI21X1
XOAI21X1_311 BUFX4_122/Y MUX2X1_28/B OAI21X1_311/C gnd NOR2X1_165/B vdd OAI21X1
XOAI21X1_388 INVX1_103/Y BUFX4_39/Y OAI21X1_388/C gnd OAI22X1_15/C vdd OAI21X1
XOAI21X1_399 INVX1_112/Y BUFX4_17/Y OAI21X1_399/C gnd INVX1_170/A vdd OAI21X1
XNAND2X1_361 BUFX4_20/Y OAI21X1_109/B gnd OAI21X1_352/C vdd NAND2X1
XNAND2X1_372 BUFX4_17/Y INVX1_94/A gnd OAI21X1_375/C vdd NAND2X1
XNAND2X1_350 BUFX4_17/Y INVX1_187/A gnd OAI21X1_339/C vdd NAND2X1
XNAND2X1_383 operand_A[41] INVX1_161/Y gnd OAI21X1_394/C vdd NAND2X1
XNAND2X1_394 INVX8_13/Y NAND2X1_394/B gnd NAND2X1_394/Y vdd NAND2X1
XFILL_7_1 gnd vdd FILL
XNAND3X1_1 NAND3X1_1/A OR2X2_45/B NOR2X1_27/Y gnd OR2X2_1/A vdd NAND3X1
XFILL_26_1_0 gnd vdd FILL
XFILL_1_1_0 gnd vdd FILL
XOAI21X1_130 MUX2X1_98/S MUX2X1_15/Y OAI21X1_130/C gnd INVX1_69/A vdd OAI21X1
XFILL_10_5_1 gnd vdd FILL
XINVX1_216 INVX1_216/A gnd INVX1_216/Y vdd INVX1
XINVX1_249 INVX1_249/A gnd INVX1_249/Y vdd INVX1
XAOI22X1_6 BUFX4_57/Y INVX2_62/Y BUFX4_6/Y AOI22X1_6/D gnd AOI22X1_6/Y vdd AOI22X1
XINVX1_205 INVX1_205/A gnd INVX1_205/Y vdd INVX1
XINVX1_238 INVX1_238/A gnd INVX1_238/Y vdd INVX1
XOAI21X1_174 AOI21X1_58/Y NOR2X1_122/B AOI21X1_60/Y gnd AOI21X1_61/C vdd OAI21X1
XOAI21X1_141 BUFX4_192/Y MUX2X1_19/Y OAI21X1_141/C gnd MUX2X1_20/B vdd OAI21X1
XINVX1_227 INVX1_227/A gnd INVX1_227/Y vdd INVX1
XOAI21X1_185 BUFX4_39/Y MUX2X1_24/Y OAI21X1_185/C gnd MUX2X1_123/A vdd OAI21X1
XOAI21X1_163 INVX1_85/Y INVX2_18/A INVX1_30/A gnd AOI21X1_54/C vdd OAI21X1
XOAI21X1_152 NOR2X1_15/Y NOR2X1_428/A NOR2X1_107/Y gnd AOI21X1_49/B vdd OAI21X1
XOAI21X1_196 INVX1_92/Y BUFX4_119/Y OAI21X1_196/C gnd INVX1_94/A vdd OAI21X1
XNAND2X1_180 MUX2X1_8/S operand_A[46] gnd OAI21X1_467/C vdd NAND2X1
XNAND2X1_49 operand_B[26] INVX2_31/Y gnd NAND2X1_50/B vdd NAND2X1
XNAND2X1_191 AND2X2_1/B NOR2X1_6/Y gnd NOR2X1_106/A vdd NAND2X1
XNAND2X1_38 operand_B[12] INVX2_21/Y gnd NAND2X1_39/B vdd NAND2X1
XNAND2X1_27 BUFX4_179/Y operand_A[4] gnd OAI21X1_12/C vdd NAND2X1
XNAND2X1_16 operand_B[17] INVX4_6/Y gnd INVX1_11/A vdd NAND2X1
XFILL_9_2_0 gnd vdd FILL
XFILL_17_1_0 gnd vdd FILL
XAOI21X1_209 INVX1_224/A OAI21X1_544/B AND2X2_33/Y gnd OAI21X1_552/B vdd AOI21X1
XAOI22X1_25 BUFX4_149/Y NOR2X1_320/B BUFX4_56/Y INVX2_82/A gnd AND2X2_39/A vdd AOI22X1
XAOI22X1_14 INVX8_17/A INVX1_182/Y INVX8_14/A INVX4_21/Y gnd NAND3X1_23/B vdd AOI22X1
XAOI22X1_58 INVX8_7/A MUX2X1_64/Y AOI22X1_58/C INVX8_9/A gnd AOI22X1_58/Y vdd AOI22X1
XAOI22X1_36 NOR2X1_25/Y BUFX4_150/Y XNOR2X1_40/Y BUFX4_140/Y gnd AOI22X1_36/Y vdd
+ AOI22X1
XAOI22X1_47 BUFX4_15/Y INVX1_272/Y AOI22X1_47/C AOI22X1_47/D gnd AOI22X1_47/Y vdd
+ AOI22X1
XOAI22X1_9 OAI22X1_9/A INVX4_23/Y OAI22X1_9/C OAI22X1_9/D gnd OAI22X1_9/Y vdd OAI22X1
XAOI21X1_91 INVX4_19/Y INVX1_144/A NOR2X1_164/Y gnd XNOR2X1_32/A vdd AOI21X1
XAOI21X1_80 NAND3X1_9/A XNOR2X1_31/Y AOI21X1_80/C gnd AOI21X1_81/B vdd AOI21X1
XNOR2X1_404 BUFX2_32/A BUFX2_31/A gnd NOR2X1_404/Y vdd NOR2X1
XNOR2X1_415 operand_A[31] INVX2_51/Y gnd NOR2X1_415/Y vdd NOR2X1
XNOR2X1_426 alu_op[1] INVX2_33/Y gnd NOR2X1_426/Y vdd NOR2X1
XNOR2X1_448 OAI21X1_10/C INVX1_302/Y gnd NOR2X1_448/Y vdd NOR2X1
XNOR2X1_459 XNOR2X1_7/Y NOR2X1_459/B gnd NOR2X1_459/Y vdd NOR2X1
XNOR2X1_437 NOR2X1_437/A NOR2X1_437/B gnd NOR2X1_437/Y vdd NOR2X1
XINVX2_29 operand_B[27] gnd INVX2_29/Y vdd INVX2
XINVX2_18 INVX2_18/A gnd INVX2_18/Y vdd INVX2
XFILL_24_4_1 gnd vdd FILL
XXOR2X1_1 operand_A[23] operand_B[23] gnd XOR2X1_1/Y vdd XOR2X1
XFILL_6_0_0 gnd vdd FILL
XFILL_7_5_1 gnd vdd FILL
XFILL_15_4_1 gnd vdd FILL
XMUX2X1_2 MUX2X1_2/A MUX2X1_2/B MUX2X1_2/S gnd MUX2X1_2/Y vdd MUX2X1
XCLKBUF1_3 clk gnd CLKBUF1_3/Y vdd CLKBUF1
XFILL_31_1 gnd vdd FILL
XNOR2X1_256 INVX2_52/Y INVX1_203/Y gnd NOR2X1_258/B vdd NOR2X1
XNOR2X1_245 OR2X2_17/B OR2X2_17/A gnd NOR2X1_245/Y vdd NOR2X1
XNOR2X1_201 operand_A[42] operand_B[42] gnd NOR2X1_202/A vdd NOR2X1
XNOR2X1_234 BUFX4_95/Y AND2X2_24/Y gnd NOR2X1_234/Y vdd NOR2X1
XBUFX4_141 NOR2X1_72/Y gnd BUFX4_141/Y vdd BUFX4
XBUFX4_174 INVX8_18/Y gnd BUFX4_174/Y vdd BUFX4
XNOR2X1_267 BUFX4_42/Y MUX2X1_45/Y gnd NOR2X1_267/Y vdd NOR2X1
XBUFX4_163 INVX8_5/Y gnd BUFX4_163/Y vdd BUFX4
XNOR2X1_212 INVX8_5/A NOR2X1_212/B gnd NOR2X1_212/Y vdd NOR2X1
XBUFX4_196 operand_B[1] gnd MUX2X1_23/S vdd BUFX4
XBUFX4_130 operand_B[2] gnd MUX2X1_99/S vdd BUFX4
XBUFX4_185 operand_B[4] gnd MUX2X1_57/S vdd BUFX4
XNOR2X1_223 MUX2X1_34/S INVX1_177/Y gnd INVX1_310/A vdd NOR2X1
XBUFX4_152 NOR2X1_89/Y gnd BUFX4_152/Y vdd BUFX4
XNOR2X1_289 BUFX4_102/Y BUFX2_56/A gnd NOR2X1_289/Y vdd NOR2X1
XNOR2X1_278 INVX1_207/A NOR2X1_278/B gnd NOR2X1_278/Y vdd NOR2X1
XOAI21X1_729 XNOR2X1_16/Y AOI21X1_51/B OAI21X1_729/C gnd NAND3X1_58/A vdd OAI21X1
XOAI21X1_718 INVX1_291/Y NOR2X1_19/B OAI21X1_718/C gnd MUX2X1_96/A vdd OAI21X1
XOAI21X1_707 INVX4_4/Y BUFX4_53/Y OAI21X1_99/C gnd OAI21X1_708/B vdd OAI21X1
XAOI21X1_392 XOR2X1_1/Y BUFX4_60/Y BUFX4_12/Y gnd NAND3X1_71/B vdd AOI21X1
XAOI21X1_381 OAI21X1_2/C OAI21X1_901/A BUFX4_96/Y gnd OAI21X1_886/C vdd AOI21X1
XINVX8_5 INVX8_5/A gnd INVX8_5/Y vdd INVX8
XAOI21X1_370 INVX8_9/A OAI21X1_870/Y OAI21X1_494/Y gnd OAI21X1_872/A vdd AOI21X1
XBUFX4_14 INVX8_19/Y gnd BUFX4_14/Y vdd BUFX4
XBUFX4_25 INVX8_2/Y gnd BUFX4_25/Y vdd BUFX4
XBUFX4_58 BUFX4_60/A gnd BUFX4_58/Y vdd BUFX4
XBUFX4_69 INVX8_1/Y gnd BUFX4_69/Y vdd BUFX4
XBUFX4_47 operand_B[0] gnd MUX2X1_5/S vdd BUFX4
XBUFX4_36 operand_B[3] gnd BUFX4_36/Y vdd BUFX4
XFILL_30_2_1 gnd vdd FILL
XOR2X2_17 OR2X2_17/A OR2X2_17/B gnd OR2X2_17/Y vdd OR2X2
XOR2X2_28 OR2X2_28/A OR2X2_28/B gnd OR2X2_28/Y vdd OR2X2
XOR2X2_39 OR2X2_39/A OR2X2_39/B gnd OR2X2_39/Y vdd OR2X2
XINVX8_17 INVX8_17/A gnd INVX8_17/Y vdd INVX8
XOAI21X1_504 BUFX4_73/Y OAI21X1_504/B OAI21X1_504/C gnd MUX2X1_51/A vdd OAI21X1
XOAI21X1_526 INVX1_210/Y BUFX4_73/Y OAI21X1_526/C gnd OAI21X1_526/Y vdd OAI21X1
XFILL_21_2_1 gnd vdd FILL
XOAI21X1_548 MUX2X1_57/S MUX2X1_52/Y OAI21X1_548/C gnd OAI21X1_548/Y vdd OAI21X1
XOAI21X1_559 OAI21X1_631/A BUFX4_37/Y OAI21X1_559/C gnd OAI21X1_560/A vdd OAI21X1
XOAI21X1_515 OAI21X1_515/A BUFX4_10/Y OAI21X1_515/C gnd OAI22X1_30/B vdd OAI21X1
XOAI21X1_537 INVX1_181/Y BUFX4_19/Y OAI21X1_537/C gnd MUX2X1_49/A vdd OAI21X1
XNAND2X1_532 NOR2X1_385/Y NOR2X1_386/Y gnd NOR2X1_389/A vdd NAND2X1
XNAND2X1_543 operand_B[54] INVX2_38/Y gnd OAI21X1_660/B vdd NAND2X1
XNAND2X1_554 operand_B[40] INVX2_47/Y gnd OAI21X1_672/B vdd NAND2X1
XNAND2X1_521 INVX1_259/Y OAI21X1_623/Y gnd NAND3X1_40/C vdd NAND2X1
XNAND2X1_510 MUX2X1_62/S OAI21X1_630/A gnd OAI21X1_593/C vdd NAND2X1
XFILL_29_3_1 gnd vdd FILL
XNAND2X1_576 BUFX4_76/Y OAI21X1_686/Y gnd OAI21X1_716/C vdd NAND2X1
XFILL_4_3_1 gnd vdd FILL
XNAND2X1_598 BUFX4_136/Y INVX1_290/A gnd OAI21X1_760/C vdd NAND2X1
XNAND2X1_565 BUFX4_37/Y OAI21X1_796/B gnd NAND3X1_56/C vdd NAND2X1
XNAND2X1_587 BUFX4_86/Y NOR2X1_142/Y gnd NAND3X1_58/C vdd NAND2X1
XFILL_12_2_1 gnd vdd FILL
XOAI21X1_323 INVX1_140/Y XOR2X1_3/A OAI21X1_323/C gnd OAI21X1_323/Y vdd OAI21X1
XOAI21X1_301 MUX2X1_30/S MUX2X1_22/Y OAI21X1_301/C gnd OAI21X1_301/Y vdd OAI21X1
XOAI21X1_312 OAI21X1_312/A BUFX4_134/Y OAI21X1_88/C gnd AND2X2_23/A vdd OAI21X1
XOAI21X1_345 NOR2X1_93/A INVX1_141/Y OAI21X1_345/C gnd OAI21X1_345/Y vdd OAI21X1
XOAI21X1_378 AND2X2_15/Y BUFX4_13/Y OAI21X1_378/C gnd OAI21X1_378/Y vdd OAI21X1
XOAI21X1_334 operand_A[38] operand_B[38] BUFX4_5/Y gnd OAI21X1_335/C vdd OAI21X1
XOAI21X1_389 OAI22X1_9/C NOR2X1_190/A AOI22X1_10/Y gnd OR2X2_18/A vdd OAI21X1
XOAI21X1_367 NOR2X1_452/B OR2X2_19/B INVX1_145/Y gnd NOR2X1_186/B vdd OAI21X1
XOAI21X1_356 NOR2X1_177/B BUFX4_41/Y INVX2_48/Y gnd OAI21X1_356/Y vdd OAI21X1
XNAND2X1_384 INVX1_169/A NOR2X1_203/Y gnd NAND2X1_384/Y vdd NAND2X1
XNAND2X1_362 INVX1_154/A INVX1_155/A gnd NAND2X1_362/Y vdd NAND2X1
XNAND2X1_395 NOR2X1_80/A MUX2X1_39/Y gnd OAI21X1_420/C vdd NAND2X1
XNAND2X1_340 AOI21X1_93/Y AOI21X1_94/Y gnd AOI21X1_95/C vdd NAND2X1
XNAND2X1_351 MUX2X1_25/S OAI21X1_339/Y gnd OAI21X1_341/C vdd NAND2X1
XNAND2X1_373 INVX8_5/A OAI21X1_375/Y gnd OAI21X1_376/C vdd NAND2X1
XOAI21X1_890 OAI21X1_890/A BUFX4_12/Y OAI21X1_890/C gnd OAI21X1_890/Y vdd OAI21X1
XFILL_7_2 gnd vdd FILL
XNAND3X1_2 INVX2_17/Y INVX1_17/Y NOR2X1_28/Y gnd OR2X2_1/B vdd NAND3X1
XFILL_26_1_1 gnd vdd FILL
XFILL_1_1_1 gnd vdd FILL
XOAI21X1_131 INVX2_53/Y BUFX4_50/Y OAI21X1_556/C gnd OAI21X1_229/B vdd OAI21X1
XOAI21X1_142 INVX2_56/Y BUFX4_48/Y OAI21X1_275/C gnd INVX1_71/A vdd OAI21X1
XOAI21X1_164 OAI21X1_164/A AOI21X1_53/Y AOI21X1_54/Y gnd AOI21X1_55/C vdd OAI21X1
XOAI21X1_120 INVX1_68/Y BUFX4_76/Y OAI21X1_120/C gnd OAI21X1_120/Y vdd OAI21X1
XOAI21X1_153 AOI21X1_49/Y AOI21X1_9/C NOR2X1_109/Y gnd AOI21X1_50/B vdd OAI21X1
XAOI22X1_7 INVX8_15/A AOI22X1_7/B AOI22X1_7/C INVX4_20/A gnd AOI22X1_7/Y vdd AOI22X1
XINVX1_239 INVX1_239/A gnd INVX1_239/Y vdd INVX1
XOAI21X1_175 INVX1_47/Y BUFX4_68/Y OAI21X1_175/C gnd OAI21X1_177/B vdd OAI21X1
XINVX1_217 INVX1_217/A gnd INVX1_217/Y vdd INVX1
XINVX1_206 INVX1_206/A gnd INVX1_206/Y vdd INVX1
XOAI21X1_197 INVX1_95/Y BUFX4_69/Y OAI21X1_197/C gnd INVX1_96/A vdd OAI21X1
XINVX1_228 INVX1_228/A gnd INVX1_228/Y vdd INVX1
XFILL_9_2_1 gnd vdd FILL
XOAI21X1_186 INVX1_86/Y BUFX4_164/Y OAI21X1_186/C gnd AND2X2_11/A vdd OAI21X1
XNAND2X1_170 BUFX4_43/Y operand_A[58] gnd OAI21X1_591/C vdd NAND2X1
XNAND2X1_192 NOR2X1_104/Y AND2X2_9/Y gnd NOR2X1_106/B vdd NAND2X1
XNAND2X1_181 NOR2X1_54/A OAI21X1_223/B gnd OAI21X1_138/C vdd NAND2X1
XNAND2X1_28 operand_A[15] INVX1_15/Y gnd INVX1_30/A vdd NAND2X1
XNAND2X1_39 NAND2X1_39/A NAND2X1_39/B gnd NAND2X1_40/B vdd NAND2X1
XNAND2X1_17 operand_A[16] INVX1_6/Y gnd NAND2X1_19/A vdd NAND2X1
XFILL_17_1_1 gnd vdd FILL
XAOI22X1_26 AOI22X1_26/A AOI22X1_26/B MUX2X1_45/Y BUFX4_42/Y gnd MUX2X1_57/B vdd AOI22X1
XAOI22X1_15 AND2X2_63/A INVX4_20/A INVX8_18/A AND2X2_64/A gnd NAND3X1_24/B vdd AOI22X1
XAOI22X1_37 BUFX4_152/Y NOR2X1_32/Y INVX2_17/Y BUFX4_60/Y gnd NAND3X1_63/B vdd AOI22X1
XAOI22X1_48 BUFX4_15/Y INVX1_271/Y NOR2X1_489/Y NAND3X1_70/Y gnd AOI22X1_48/Y vdd
+ AOI22X1
XAOI21X1_70 NOR2X1_137/Y INVX4_16/A NOR2X1_138/Y gnd AOI21X1_70/Y vdd AOI21X1
XAOI21X1_81 AOI21X1_81/A AOI21X1_81/B NOR2X1_152/Y gnd AOI21X1_81/Y vdd AOI21X1
XAOI21X1_92 BUFX4_36/Y AND2X2_23/A INVX1_135/A gnd INVX1_221/A vdd AOI21X1
XNOR2X1_416 operand_A[59] INVX1_242/Y gnd NOR2X1_416/Y vdd NOR2X1
XNOR2X1_405 BUFX2_28/A BUFX2_27/A gnd NOR2X1_405/Y vdd NOR2X1
XNOR2X1_438 NOR2X1_438/A NOR2X1_438/B gnd NOR2X1_438/Y vdd NOR2X1
XNOR2X1_427 BUFX4_179/Y NAND3X1_7/Y gnd NOR2X1_427/Y vdd NOR2X1
XNOR2X1_449 MUX2X1_32/S NOR2X1_449/B gnd NOR2X1_450/B vdd NOR2X1
XINVX2_19 INVX2_19/A gnd INVX2_19/Y vdd INVX2
XFILL_6_0_1 gnd vdd FILL
XXOR2X1_2 operand_B[19] operand_A[19] gnd XOR2X1_2/Y vdd XOR2X1
XMUX2X1_3 operand_A[13] operand_A[14] MUX2X1_3/S gnd MUX2X1_3/Y vdd MUX2X1
XCLKBUF1_4 clk gnd CLKBUF1_4/Y vdd CLKBUF1
XBUFX4_120 INVX8_3/Y gnd BUFX4_120/Y vdd BUFX4
XNOR2X1_246 BUFX4_32/Y AND2X2_26/Y gnd NOR2X1_246/Y vdd NOR2X1
XNOR2X1_257 operand_A[49] operand_B[49] gnd NOR2X1_258/A vdd NOR2X1
XNOR2X1_279 INVX2_78/Y INVX1_216/A gnd NOR2X1_286/B vdd NOR2X1
XNOR2X1_202 NOR2X1_202/A NOR2X1_202/B gnd INVX1_169/A vdd NOR2X1
XBUFX4_153 NOR2X1_89/Y gnd BUFX4_153/Y vdd BUFX4
XFILL_24_1 gnd vdd FILL
XBUFX4_142 NOR2X1_72/Y gnd NAND3X1_9/A vdd BUFX4
XNOR2X1_224 OR2X2_8/B NOR2X1_224/B gnd NOR2X1_224/Y vdd NOR2X1
XBUFX4_175 INVX8_18/Y gnd OR2X2_25/B vdd BUFX4
XNOR2X1_235 OR2X2_43/B OAI21X1_74/Y gnd NOR2X1_235/Y vdd NOR2X1
XNOR2X1_268 INVX8_15/Y NOR2X1_268/B gnd OR2X2_31/A vdd NOR2X1
XBUFX4_131 operand_B[2] gnd BUFX4_131/Y vdd BUFX4
XNOR2X1_213 OR2X2_43/B OAI22X1_19/A gnd NOR2X1_213/Y vdd NOR2X1
XBUFX4_186 operand_B[4] gnd BUFX4_186/Y vdd BUFX4
XBUFX4_164 INVX8_5/Y gnd BUFX4_164/Y vdd BUFX4
XOAI21X1_719 INVX1_286/Y BUFX4_74/Y OAI21X1_719/C gnd MUX2X1_110/A vdd OAI21X1
XOAI21X1_708 BUFX4_192/Y OAI21X1_708/B OAI21X1_708/C gnd OAI21X1_708/Y vdd OAI21X1
XINVX8_6 INVX8_6/A gnd INVX8_6/Y vdd INVX8
XAOI21X1_393 INVX8_6/A XNOR2X1_46/Y NAND3X1_71/Y gnd AOI22X1_54/C vdd AOI21X1
XAOI21X1_371 BUFX4_91/Y AOI22X1_19/B OAI21X1_871/Y gnd OAI21X1_872/B vdd AOI21X1
XAOI21X1_382 BUFX4_163/Y MUX2X1_107/B INVX8_4/A gnd OAI21X1_887/C vdd AOI21X1
XAOI21X1_360 XNOR2X1_22/Y NOR2X1_476/Y BUFX4_31/Y gnd OAI21X1_857/C vdd AOI21X1
XBUFX4_59 BUFX4_60/A gnd INVX8_14/A vdd BUFX4
XBUFX4_48 operand_B[0] gnd BUFX4_48/Y vdd BUFX4
XBUFX4_37 operand_B[3] gnd BUFX4_37/Y vdd BUFX4
XBUFX4_26 INVX8_2/Y gnd OR2X2_39/B vdd BUFX4
XBUFX4_15 INVX8_19/Y gnd BUFX4_15/Y vdd BUFX4
XOR2X2_29 OR2X2_29/A OR2X2_29/B gnd OR2X2_29/Y vdd OR2X2
XOR2X2_18 OR2X2_18/A OR2X2_8/B gnd OR2X2_18/Y vdd OR2X2
XINVX8_18 INVX8_18/A gnd INVX8_18/Y vdd INVX8
XOAI21X1_505 NOR2X1_267/Y NOR2X1_266/Y MUX2X1_49/S gnd OAI21X1_506/C vdd OAI21X1
XOAI21X1_527 INVX1_217/Y MUX2X1_66/S OAI21X1_527/C gnd MUX2X1_61/A vdd OAI21X1
XOAI21X1_538 NOR2X1_493/B BUFX4_10/Y OAI21X1_538/C gnd OAI21X1_539/A vdd OAI21X1
XOAI21X1_549 INVX1_147/A INVX8_5/A OAI21X1_549/C gnd NOR2X1_294/B vdd OAI21X1
XOAI21X1_516 OAI22X1_30/B NOR2X1_274/Y BUFX4_78/Y gnd OAI21X1_516/Y vdd OAI21X1
XNAND2X1_533 NOR2X1_387/Y NOR2X1_388/Y gnd NOR2X1_389/B vdd NAND2X1
XNAND2X1_544 operand_B[53] INVX2_53/Y gnd OAI21X1_661/C vdd NAND2X1
XNAND2X1_511 INVX1_239/A NOR2X1_345/Y gnd INVX1_247/A vdd NAND2X1
XNAND2X1_555 NOR2X1_218/Y OAI21X1_672/Y gnd NAND2X1_555/Y vdd NAND2X1
XNAND2X1_522 MUX2X1_8/S operand_A[61] gnd OAI21X1_624/C vdd NAND2X1
XNAND2X1_588 INVX8_1/A MUX2X1_77/Y gnd OAI21X1_733/C vdd NAND2X1
XNAND2X1_500 BUFX4_70/Y INVX1_238/Y gnd OAI21X1_577/C vdd NAND2X1
XNAND2X1_577 BUFX4_74/Y OAI21X1_683/Y gnd OAI21X1_717/C vdd NAND2X1
XNAND2X1_566 BUFX4_116/Y AND2X2_11/A gnd OAI21X1_695/C vdd NAND2X1
XNAND2X1_599 MUX2X1_27/S OAI21X1_703/Y gnd OAI21X1_761/C vdd NAND2X1
XAOI21X1_190 AOI21X1_190/A OAI21X1_509/Y NOR2X1_275/Y gnd DFFPOSX1_52/D vdd AOI21X1
XFILL_31_5_0 gnd vdd FILL
XOAI21X1_346 INVX2_66/Y INVX2_67/Y OAI21X1_346/C gnd OAI21X1_347/B vdd OAI21X1
XOAI21X1_335 OAI22X1_9/A OR2X2_12/B OAI21X1_335/C gnd NOR2X1_171/A vdd OAI21X1
XFILL_22_5_0 gnd vdd FILL
XOAI21X1_302 BUFX4_16/Y NOR2X1_222/B OAI21X1_302/C gnd INVX1_133/A vdd OAI21X1
XOAI21X1_324 INVX1_106/Y BUFX4_122/Y OAI21X1_324/C gnd OAI21X1_443/B vdd OAI21X1
XOAI21X1_313 INVX1_221/A BUFX4_164/Y OAI21X1_313/C gnd AND2X2_56/A vdd OAI21X1
XOAI21X1_357 INVX1_148/A INVX1_143/A NOR2X1_174/A gnd OAI21X1_357/Y vdd OAI21X1
XOAI21X1_379 INVX1_162/Y OAI21X1_379/B OAI21X1_379/C gnd OAI21X1_379/Y vdd OAI21X1
XOAI21X1_368 INVX1_98/Y XOR2X1_7/A XOR2X1_4/A gnd OAI21X1_369/C vdd OAI21X1
XNAND2X1_341 operand_A[38] operand_B[38] gnd INVX1_143/A vdd NAND2X1
XNAND2X1_363 OR2X2_12/B INVX1_148/A gnd NOR2X1_183/B vdd NAND2X1
XNAND2X1_374 INVX8_18/A AND2X2_57/A gnd NAND3X1_17/C vdd NAND2X1
XNAND2X1_396 OAI21X1_419/Y OAI21X1_420/C gnd AOI22X1_12/A vdd NAND2X1
XNAND2X1_330 BUFX4_162/Y NOR2X1_166/Y gnd NOR2X1_444/B vdd NAND2X1
XNAND2X1_385 BUFX4_17/Y INVX1_114/A gnd OAI21X1_399/C vdd NAND2X1
XNAND2X1_352 BUFX4_17/Y OAI21X1_50/B gnd OAI21X1_340/C vdd NAND2X1
XFILL_13_5_0 gnd vdd FILL
XOAI21X1_891 OAI21X1_901/A OAI21X1_2/C NAND2X1_8/A gnd AND2X2_71/A vdd OAI21X1
XOAI21X1_880 XOR2X1_2/Y OAI21X1_880/B OAI21X1_880/C gnd AOI22X1_49/D vdd OAI21X1
XNAND3X1_3 AND2X2_4/Y NAND3X1_3/B OAI22X1_2/Y gnd NOR2X1_91/B vdd NAND3X1
XINVX1_207 INVX1_207/A gnd INVX1_207/Y vdd INVX1
XOAI21X1_165 operand_A[31] INVX2_51/Y NOR2X1_97/A gnd OAI21X1_166/C vdd OAI21X1
XAOI22X1_8 BUFX4_58/Y INVX2_65/Y BUFX4_5/Y OR2X2_11/Y gnd AOI22X1_8/Y vdd AOI22X1
XOAI21X1_198 INVX2_45/Y MUX2X1_3/S OAI21X1_198/C gnd INVX1_97/A vdd OAI21X1
XOAI21X1_154 AOI21X1_50/Y AOI21X1_47/C AOI22X1_4/C gnd INVX1_78/A vdd OAI21X1
XOAI21X1_143 INVX2_50/Y BUFX4_50/Y OAI21X1_217/C gnd OAI21X1_703/B vdd OAI21X1
XOAI21X1_176 NOR2X1_82/A INVX1_49/A OAI21X1_176/C gnd OAI21X1_176/Y vdd OAI21X1
XOAI21X1_132 MUX2X1_23/S MUX2X1_16/Y OAI21X1_132/C gnd MUX2X1_30/A vdd OAI21X1
XOAI21X1_187 BUFX4_190/Y OAI21X1_55/Y OAI21X1_187/C gnd OAI21X1_187/Y vdd OAI21X1
XOAI21X1_121 INVX1_67/Y MUX2X1_2/S OAI21X1_121/C gnd INVX1_149/A vdd OAI21X1
XOAI21X1_110 INVX2_9/Y MUX2X1_7/S INVX2_10/A gnd INVX1_101/A vdd OAI21X1
XINVX1_218 operand_B[53] gnd INVX1_218/Y vdd INVX1
XINVX1_229 INVX1_229/A gnd INVX1_229/Y vdd INVX1
XNAND2X1_193 operand_B[30] INVX2_35/Y gnd INVX1_76/A vdd NAND2X1
XNAND2X1_171 BUFX4_191/Y OAI21X1_126/Y gnd OAI21X1_127/C vdd NAND2X1
XNAND2X1_182 BUFX4_134/Y OAI21X1_265/B gnd OAI21X1_139/C vdd NAND2X1
XNAND2X1_29 operand_B[15] INVX2_15/Y gnd INVX1_85/A vdd NAND2X1
XNAND2X1_160 BUFX4_46/Y operand_A[8] gnd OAI21X1_116/C vdd NAND2X1
XNAND2X1_18 operand_B[16] INVX2_6/Y gnd NAND2X1_19/B vdd NAND2X1
XAOI22X1_27 BUFX4_56/Y OR2X2_34/B BUFX4_4/Y INVX1_244/Y gnd AOI22X1_27/Y vdd AOI22X1
XAOI22X1_16 INVX8_17/A NOR2X1_231/B BUFX4_57/Y INVX1_186/A gnd AOI22X1_16/Y vdd AOI22X1
XAOI22X1_38 AOI22X1_38/A BUFX4_90/Y INVX8_10/A AOI22X1_38/D gnd AND2X2_58/A vdd AOI22X1
XAOI22X1_49 BUFX4_15/Y INVX1_270/Y AOI22X1_49/C AOI22X1_49/D gnd AOI22X1_49/Y vdd
+ AOI22X1
XFILL_27_4_0 gnd vdd FILL
XFILL_2_4_0 gnd vdd FILL
XAOI21X1_82 INVX1_108/A NOR2X1_155/Y AOI21X1_82/C gnd AOI21X1_82/Y vdd AOI21X1
XAOI21X1_60 AOI21X1_60/A NOR2X1_121/Y AOI21X1_60/C gnd AOI21X1_60/Y vdd AOI21X1
XAOI21X1_71 BUFX4_136/Y NOR2X1_139/Y INVX1_109/A gnd AOI21X1_71/Y vdd AOI21X1
XAOI21X1_93 INVX4_20/A AND2X2_56/A AOI21X1_93/C gnd AOI21X1_93/Y vdd AOI21X1
XFILL_10_3_0 gnd vdd FILL
XNOR2X1_417 operand_A[58] INVX2_83/Y gnd NOR2X1_417/Y vdd NOR2X1
XNOR2X1_406 NOR2X1_406/A NOR2X1_406/B gnd NOR2X1_406/Y vdd NOR2X1
XFILL_18_4_0 gnd vdd FILL
XNOR2X1_428 NOR2X1_428/A BUFX4_27/Y gnd NOR2X1_428/Y vdd NOR2X1
XNOR2X1_439 NOR2X1_439/A INVX1_297/Y gnd NOR2X1_441/A vdd NOR2X1
XXOR2X1_3 XOR2X1_3/A operand_A[1] gnd XOR2X1_3/Y vdd XOR2X1
XMUX2X1_4 operand_A[9] operand_A[10] MUX2X1_4/S gnd MUX2X1_4/Y vdd MUX2X1
XCLKBUF1_5 clk gnd CLKBUF1_5/Y vdd CLKBUF1
XBUFX4_143 NOR2X1_72/Y gnd BUFX4_143/Y vdd BUFX4
XBUFX4_121 INVX8_3/Y gnd MUX2X1_66/S vdd BUFX4
XBUFX4_132 operand_B[2] gnd MUX2X1_51/S vdd BUFX4
XBUFX4_110 operand_B[5] gnd INVX8_4/A vdd BUFX4
XBUFX4_154 INVX8_14/Y gnd BUFX4_154/Y vdd BUFX4
XNOR2X1_236 BUFX4_101/Y BUFX2_49/A gnd NOR2X1_236/Y vdd NOR2X1
XNOR2X1_214 BUFX4_102/Y BUFX2_46/A gnd NOR2X1_214/Y vdd NOR2X1
XNOR2X1_258 NOR2X1_258/A NOR2X1_258/B gnd INVX1_204/A vdd NOR2X1
XNOR2X1_269 operand_A[51] operand_B[51] gnd INVX1_214/A vdd NOR2X1
XNOR2X1_203 NOR2X1_203/A AND2X2_17/Y gnd NOR2X1_203/Y vdd NOR2X1
XNOR2X1_247 OR2X2_29/Y NOR2X1_247/B gnd INVX1_200/A vdd NOR2X1
XNOR2X1_225 BUFX4_99/Y BUFX2_48/A gnd NOR2X1_225/Y vdd NOR2X1
XFILL_17_1 gnd vdd FILL
XBUFX4_176 INVX8_18/Y gnd OR2X2_16/B vdd BUFX4
XBUFX4_187 operand_B[1] gnd INVX8_1/A vdd BUFX4
XBUFX4_165 INVX8_5/Y gnd MUX2X1_64/S vdd BUFX4
XOAI21X1_709 INVX4_6/Y MUX2X1_8/S OAI21X1_96/C gnd OAI21X1_710/B vdd OAI21X1
XFILL_24_2_0 gnd vdd FILL
XINVX8_7 INVX8_7/A gnd INVX8_7/Y vdd INVX8
XAOI21X1_361 XNOR2X1_22/Y OAI21X1_859/A OAI21X1_859/Y gnd NOR2X1_479/A vdd AOI21X1
XAOI21X1_350 NAND3X1_65/Y AOI21X1_350/B NOR2X1_469/Y gnd DFFPOSX1_14/D vdd AOI21X1
XDFFPOSX1_60 BUFX2_62/A CLKBUF1_5/Y DFFPOSX1_60/D gnd vdd DFFPOSX1
XAOI21X1_394 XNOR2X1_29/Y OAI21X1_23/A BUFX4_31/Y gnd OAI21X1_909/C vdd AOI21X1
XAOI21X1_383 INVX8_12/A OAI21X1_523/Y OAI21X1_888/Y gnd OAI21X1_889/A vdd AOI21X1
XAOI21X1_372 INVX4_26/Y INVX8_14/A BUFX4_12/Y gnd AND2X2_70/B vdd AOI21X1
XBUFX4_27 INVX8_6/Y gnd BUFX4_27/Y vdd BUFX4
XBUFX4_16 INVX8_2/Y gnd BUFX4_16/Y vdd BUFX4
XBUFX4_49 operand_B[0] gnd MUX2X1_1/S vdd BUFX4
XBUFX4_38 operand_B[3] gnd BUFX4_38/Y vdd BUFX4
XFILL_7_3_0 gnd vdd FILL
XFILL_15_2_0 gnd vdd FILL
XOR2X2_19 OR2X2_19/A OR2X2_19/B gnd OR2X2_19/Y vdd OR2X2
XOAI21X1_517 NOR2X1_273/A NOR2X1_271/B INVX1_214/Y gnd OAI21X1_518/C vdd OAI21X1
XOAI21X1_528 OR2X2_7/B MUX2X1_47/Y OAI21X1_528/C gnd MUX2X1_48/A vdd OAI21X1
XOAI21X1_539 OAI21X1_539/A NOR2X1_287/Y BUFX4_79/Y gnd NAND3X1_32/C vdd OAI21X1
XOAI21X1_506 OAI21X1_506/A MUX2X1_49/S OAI21X1_506/C gnd NOR2X1_268/B vdd OAI21X1
XINVX8_19 OR2X2_48/A gnd INVX8_19/Y vdd INVX8
XNAND2X1_534 NOR2X1_391/Y NOR2X1_392/Y gnd NOR2X1_393/B vdd NAND2X1
XNAND2X1_545 operand_B[52] INVX2_40/Y gnd OAI21X1_661/B vdd NAND2X1
XNAND2X1_512 INVX1_237/A INVX1_249/A gnd INVX1_248/A vdd NAND2X1
XNAND2X1_523 INVX8_13/Y NAND2X1_523/B gnd NAND2X1_523/Y vdd NAND2X1
XNAND2X1_556 alu_op[3] INVX1_43/Y gnd NAND2X1_556/Y vdd NAND2X1
XNAND2X1_589 INVX8_3/A MUX2X1_20/A gnd OAI21X1_734/C vdd NAND2X1
XNAND2X1_501 MUX2X1_87/S OAI21X1_535/Y gnd OAI21X1_578/C vdd NAND2X1
XNAND2X1_578 BUFX4_125/Y MUX2X1_110/B gnd OAI21X1_718/C vdd NAND2X1
XNAND2X1_567 OAI21X1_700/Y NAND2X1_567/B gnd NAND2X1_567/Y vdd NAND2X1
XAOI21X1_191 NOR2X1_278/Y AND2X2_26/A OAI21X1_518/Y gnd INVX1_216/A vdd AOI21X1
XAOI21X1_180 BUFX4_159/Y OAI21X1_250/Y INVX4_11/A gnd NOR2X1_487/B vdd AOI21X1
XFILL_31_5_1 gnd vdd FILL
XFILL_30_0_0 gnd vdd FILL
XOAI21X1_347 INVX1_148/Y OAI21X1_347/B OAI21X1_347/C gnd OAI21X1_347/Y vdd OAI21X1
XOAI21X1_358 AOI21X1_82/Y OR2X2_17/B OAI21X1_358/C gnd INVX1_153/A vdd OAI21X1
XOAI21X1_336 INVX2_66/Y MUX2X1_1/S OAI21X1_75/C gnd INVX1_159/A vdd OAI21X1
XFILL_22_5_1 gnd vdd FILL
XFILL_21_0_0 gnd vdd FILL
XOAI21X1_303 AOI21X1_86/Y BUFX4_159/Y OAI21X1_304/C gnd AND2X2_55/A vdd OAI21X1
XOAI21X1_314 INVX1_101/Y MUX2X1_23/S MUX2X1_87/S gnd OAI21X1_315/C vdd OAI21X1
XOAI21X1_369 OAI21X1_369/A BUFX4_35/Y OAI21X1_369/C gnd OR2X2_43/A vdd OAI21X1
XOAI21X1_325 INVX1_139/Y BUFX4_23/Y OAI21X1_325/C gnd MUX2X1_49/B vdd OAI21X1
XNAND2X1_320 BUFX4_16/Y OAI21X1_301/Y gnd OAI21X1_302/C vdd NAND2X1
XBUFX4_1 BUFX4_6/A gnd BUFX4_1/Y vdd BUFX4
XNAND2X1_342 INVX2_66/Y INVX2_67/Y gnd NAND2X1_343/B vdd NAND2X1
XNAND2X1_353 operand_A[39] operand_B[39] gnd NOR2X1_174/A vdd NAND2X1
XNAND2X1_375 BUFX2_43/A BUFX4_13/Y gnd OAI21X1_378/C vdd NAND2X1
XFILL_29_1_0 gnd vdd FILL
XNAND2X1_364 INVX1_157/A INVX1_127/A gnd INVX1_158/A vdd NAND2X1
XNAND2X1_386 BUFX4_75/Y INVX1_171/Y gnd OAI21X1_401/C vdd NAND2X1
XNAND2X1_397 BUFX4_21/Y OAI21X1_268/Y gnd OAI22X1_18/B vdd NAND2X1
XNAND2X1_331 BUFX4_122/Y MUX2X1_28/A gnd NOR2X1_228/B vdd NAND2X1
XFILL_4_1_0 gnd vdd FILL
XINVX4_1 INVX4_1/A gnd INVX4_1/Y vdd INVX4
XFILL_13_5_1 gnd vdd FILL
XFILL_12_0_0 gnd vdd FILL
XOAI21X1_892 AND2X2_71/A AND2X2_71/B BUFX4_140/Y gnd OAI21X1_898/B vdd OAI21X1
XOAI21X1_870 AND2X2_69/Y OAI21X1_870/B BUFX4_77/Y gnd OAI21X1_870/Y vdd OAI21X1
XOAI21X1_881 NOR2X1_486/Y OR2X2_47/B NAND2X1_9/Y gnd XNOR2X1_43/A vdd OAI21X1
XNAND3X1_4 NAND3X1_4/A NAND3X1_4/B NAND3X1_4/C gnd NAND3X1_4/Y vdd NAND3X1
XAOI22X1_9 BUFX4_153/Y INVX1_143/Y OR2X2_12/Y AOI22X1_9/D gnd AOI22X1_9/Y vdd AOI22X1
XINVX1_208 INVX1_208/A gnd INVX1_208/Y vdd INVX1
XINVX1_219 INVX1_219/A gnd INVX1_219/Y vdd INVX1
XOAI21X1_166 INVX2_50/Y operand_B[31] OAI21X1_166/C gnd AOI21X1_56/C vdd OAI21X1
XOAI21X1_155 AOI22X1_4/C INVX1_77/Y NOR2X1_111/Y gnd AOI21X1_65/A vdd OAI21X1
XOAI21X1_144 INVX1_71/Y BUFX4_72/Y OAI21X1_144/C gnd MUX2X1_20/A vdd OAI21X1
XOAI21X1_199 INVX1_97/Y MUX2X1_98/S OAI21X1_199/C gnd OAI21X1_199/Y vdd OAI21X1
XOAI21X1_177 MUX2X1_30/S OAI21X1_177/B OAI21X1_177/C gnd OAI21X1_365/B vdd OAI21X1
XOAI21X1_133 INVX1_69/Y BUFX4_133/Y OAI21X1_133/C gnd MUX2X1_36/B vdd OAI21X1
XOAI21X1_111 INVX2_11/Y MUX2X1_3/S OAI21X1_111/C gnd INVX1_65/A vdd OAI21X1
XOAI21X1_188 BUFX4_192/Y INVX1_36/A OAI21X1_188/C gnd INVX1_89/A vdd OAI21X1
XOAI21X1_100 INVX1_60/Y BUFX4_67/Y OAI21X1_100/C gnd OAI21X1_100/Y vdd OAI21X1
XOAI21X1_122 INVX1_66/Y OR2X2_39/B OAI21X1_122/C gnd OAI21X1_123/A vdd OAI21X1
XNAND2X1_150 BUFX4_48/Y operand_A[28] gnd OAI21X1_105/C vdd NAND2X1
XNAND2X1_161 NOR2X1_54/A OAI21X1_211/B gnd OAI21X1_117/C vdd NAND2X1
XNAND2X1_19 NAND2X1_19/A NAND2X1_19/B gnd OAI21X1_7/C vdd NAND2X1
XNAND2X1_183 MUX2X1_9/S operand_A[38] gnd OAI21X1_348/C vdd NAND2X1
XNAND2X1_172 XOR2X1_4/A NOR2X1_177/B gnd OAI21X1_134/C vdd NAND2X1
XNAND2X1_194 operand_A[1] BUFX4_66/Y gnd AOI21X1_48/A vdd NAND2X1
XAOI22X1_28 BUFX4_149/Y INVX1_257/A BUFX4_4/Y INVX1_255/Y gnd AOI22X1_28/Y vdd AOI22X1
XAOI22X1_17 INVX8_17/A INVX1_194/Y BUFX4_58/Y INVX4_22/Y gnd NAND3X1_28/B vdd AOI22X1
XAOI22X1_39 BUFX4_11/Y INVX1_264/Y AND2X2_58/Y AOI22X1_39/D gnd AOI22X1_39/Y vdd AOI22X1
XFILL_5_1 gnd vdd FILL
XBUFX2_60 OR2X2_37/B gnd result[57] vdd BUFX2
XFILL_27_4_1 gnd vdd FILL
XFILL_2_4_1 gnd vdd FILL
XFILL_10_3_1 gnd vdd FILL
XAOI21X1_83 INVX4_19/Y INVX2_64/Y AOI21X1_83/C gnd AOI21X1_83/Y vdd AOI21X1
XAOI21X1_61 NOR2X1_122/Y OAI21X1_32/Y AOI21X1_61/C gnd AOI21X1_62/B vdd AOI21X1
XAOI21X1_50 OAI21X1_19/C AOI21X1_50/B AOI21X1_50/C gnd AOI21X1_50/Y vdd AOI21X1
XOAI21X1_1 INVX1_3/Y NOR2X1_4/Y XOR2X1_1/Y gnd NOR2X1_6/B vdd OAI21X1
XAOI21X1_72 AOI21X1_72/A AOI21X1_72/B BUFX4_7/Y gnd AOI21X1_75/B vdd AOI21X1
XAOI21X1_94 BUFX4_86/Y AOI21X1_94/B NOR2X1_168/Y gnd AOI21X1_94/Y vdd AOI21X1
XFILL_9_0_0 gnd vdd FILL
XNOR2X1_407 NOR2X1_407/A NOR2X1_407/B gnd AND2X2_45/B vdd NOR2X1
XNOR2X1_418 operand_A[39] INVX2_70/Y gnd NOR2X1_418/Y vdd NOR2X1
XFILL_18_4_1 gnd vdd FILL
XNOR2X1_429 BUFX4_14/Y NOR2X1_429/B gnd NOR2X1_429/Y vdd NOR2X1
XMUX2X1_5 operand_A[61] operand_A[60] MUX2X1_5/S gnd MUX2X1_5/Y vdd MUX2X1
XXOR2X1_4 XOR2X1_4/A operand_A[3] gnd XOR2X1_4/Y vdd XOR2X1
XCLKBUF1_6 clk gnd DFFSR_1/CLK vdd CLKBUF1
XNOR2X1_215 BUFX4_101/Y BUFX2_47/A gnd NOR2X1_215/Y vdd NOR2X1
XBUFX4_144 INVX8_16/Y gnd OAI22X1_7/C vdd BUFX4
XNOR2X1_204 BUFX4_163/Y INVX1_170/Y gnd NOR2X1_204/Y vdd NOR2X1
XBUFX4_166 INVX8_5/Y gnd MUX2X1_49/S vdd BUFX4
XBUFX4_122 INVX8_3/Y gnd BUFX4_122/Y vdd BUFX4
XBUFX4_188 operand_B[1] gnd XOR2X1_3/A vdd BUFX4
XBUFX4_133 operand_B[2] gnd BUFX4_133/Y vdd BUFX4
XBUFX4_111 operand_B[5] gnd BUFX4_111/Y vdd BUFX4
XBUFX4_177 operand_B[4] gnd INVX8_5/A vdd BUFX4
XBUFX4_155 INVX8_14/Y gnd BUFX4_155/Y vdd BUFX4
XBUFX4_100 DFFSR_1/Q gnd BUFX4_100/Y vdd BUFX4
XNOR2X1_259 INVX1_201/A AND2X2_26/Y gnd NOR2X1_259/Y vdd NOR2X1
XNOR2X1_237 BUFX4_101/Y BUFX2_50/A gnd NOR2X1_237/Y vdd NOR2X1
XNOR2X1_248 OR2X2_29/Y NOR2X1_248/B gnd NOR2X1_251/B vdd NOR2X1
XNOR2X1_226 AND2X2_21/Y NOR2X1_226/B gnd NOR2X1_226/Y vdd NOR2X1
XFILL_17_2 gnd vdd FILL
XFILL_24_2_1 gnd vdd FILL
XAOI21X1_395 NAND2X1_59/B OAI21X1_34/A OAI21X1_910/Y gnd NOR2X1_499/A vdd AOI21X1
XAOI21X1_384 BUFX4_108/Y XNOR2X1_44/Y NAND2X1_634/Y gnd OAI21X1_890/A vdd AOI21X1
XAOI21X1_362 INVX8_5/A MUX2X1_21/B OAI21X1_860/Y gnd OAI21X1_862/B vdd AOI21X1
XAOI21X1_351 NOR2X1_27/Y OAI21X1_833/A INVX1_312/Y gnd NOR2X1_472/B vdd AOI21X1
XAOI21X1_340 NOR2X1_34/Y BUFX4_152/Y BUFX4_11/Y gnd NAND2X1_618/A vdd AOI21X1
XINVX8_8 INVX8_8/A gnd INVX8_8/Y vdd INVX8
XAOI21X1_373 BUFX4_138/Y XNOR2X1_42/Y OAI21X1_872/Y gnd AOI22X1_47/C vdd AOI21X1
XDFFPOSX1_50 BUFX2_52/A CLKBUF1_4/Y DFFPOSX1_50/D gnd vdd DFFPOSX1
XDFFPOSX1_61 BUFX2_63/A CLKBUF1_5/Y DFFPOSX1_61/D gnd vdd DFFPOSX1
XBUFX4_28 INVX8_6/Y gnd BUFX4_28/Y vdd BUFX4
XBUFX4_39 operand_B[3] gnd BUFX4_39/Y vdd BUFX4
XFILL_7_3_1 gnd vdd FILL
XBUFX4_17 INVX8_2/Y gnd BUFX4_17/Y vdd BUFX4
XFILL_15_2_1 gnd vdd FILL
XOAI21X1_529 NAND3X1_31/Y OAI21X1_529/B BUFX4_102/Y gnd OAI21X1_530/C vdd OAI21X1
XOAI21X1_518 INVX1_208/A NOR2X1_278/B OAI21X1_518/C gnd OAI21X1_518/Y vdd OAI21X1
XOAI21X1_507 OAI21X1_875/A OR2X2_16/B AND2X2_31/Y gnd OR2X2_31/B vdd OAI21X1
XNAND2X1_502 NOR2X1_80/A NOR2X1_197/Y gnd OAI21X1_917/A vdd NAND2X1
XNAND2X1_546 operand_B[37] INVX2_55/Y gnd OAI21X1_664/C vdd NAND2X1
XNAND2X1_568 BUFX4_72/Y MUX2X1_77/Y gnd OAI21X1_703/C vdd NAND2X1
XNAND2X1_524 NAND2X1_524/A OAI22X1_21/Y gnd NAND2X1_524/Y vdd NAND2X1
XNAND2X1_557 BUFX4_190/Y OAI21X1_676/Y gnd OAI21X1_677/C vdd NAND2X1
XNAND2X1_513 INVX8_5/A MUX2X1_40/Y gnd NAND2X1_513/Y vdd NAND2X1
XNAND2X1_579 BUFX4_74/Y MUX2X1_76/B gnd OAI21X1_719/C vdd NAND2X1
XNAND2X1_535 NOR2X1_397/Y NOR2X1_400/Y gnd NOR2X1_407/A vdd NAND2X1
XAOI21X1_170 OAI21X1_473/Y AND2X2_28/Y NOR2X1_240/Y gnd DFFPOSX1_49/D vdd AOI21X1
XAOI21X1_192 NOR2X1_281/Y OAI21X1_501/Y OAI21X1_520/Y gnd NOR2X1_312/B vdd AOI21X1
XAOI21X1_181 MUX2X1_64/S OAI21X1_261/B OAI21X1_502/Y gnd OAI22X1_29/D vdd AOI21X1
XFILL_30_0_1 gnd vdd FILL
XOAI21X1_359 INVX1_77/A OR2X2_17/Y INVX1_153/Y gnd INVX1_155/A vdd OAI21X1
XOAI21X1_348 INVX2_69/Y BUFX4_50/Y OAI21X1_348/C gnd OAI21X1_348/Y vdd OAI21X1
XFILL_21_0_1 gnd vdd FILL
XOAI21X1_337 INVX1_130/Y BUFX4_75/Y OAI21X1_337/C gnd OAI21X1_337/Y vdd OAI21X1
XOAI21X1_304 INVX1_133/Y BUFX4_159/Y OAI21X1_304/C gnd INVX1_296/A vdd OAI21X1
XOAI21X1_315 OAI21X1_315/A BUFX4_136/Y OAI21X1_315/C gnd NOR2X1_166/B vdd OAI21X1
XOAI21X1_326 INVX1_138/Y MUX2X1_25/S OAI21X1_326/C gnd AOI21X1_94/B vdd OAI21X1
XNAND2X1_343 INVX1_143/A NAND2X1_343/B gnd OR2X2_12/B vdd NAND2X1
XNAND2X1_354 INVX2_69/Y INVX2_70/Y gnd NAND2X1_355/B vdd NAND2X1
XNAND2X1_321 MUX2X1_30/S MUX2X1_23/Y gnd NOR2X1_222/B vdd NAND2X1
XNAND2X1_310 BUFX4_120/Y INVX1_96/A gnd OAI21X1_292/C vdd NAND2X1
XNAND2X1_332 MUX2X1_27/S OAI21X1_215/Y gnd OAI21X1_319/C vdd NAND2X1
XBUFX4_2 BUFX4_6/A gnd BUFX4_2/Y vdd BUFX4
XFILL_29_1_1 gnd vdd FILL
XNAND2X1_376 operand_A[40] INVX1_152/Y gnd AND2X2_16/B vdd NAND2X1
XNAND2X1_398 operand_B[43] INVX2_73/Y gnd NAND3X1_21/C vdd NAND2X1
XNAND2X1_387 MUX2X1_51/S OAI21X1_337/Y gnd OAI21X1_402/C vdd NAND2X1
XNAND2X1_365 BUFX4_25/Y OAI21X1_178/Y gnd NOR2X1_317/B vdd NAND2X1
XFILL_4_1_1 gnd vdd FILL
XINVX4_2 operand_A[28] gnd INVX4_2/Y vdd INVX4
XFILL_12_0_1 gnd vdd FILL
XOAI21X1_893 XNOR2X1_44/A XNOR2X1_13/Y INVX1_321/A gnd XNOR2X1_45/A vdd OAI21X1
XOAI21X1_871 OAI21X1_871/A BUFX4_172/Y BUFX4_116/Y gnd OAI21X1_871/Y vdd OAI21X1
XOAI21X1_882 INVX1_318/Y NOR2X1_75/A OAI21X1_882/C gnd OAI21X1_882/Y vdd OAI21X1
XOAI21X1_860 MUX2X1_122/Y BUFX4_186/Y BUFX4_78/Y gnd OAI21X1_860/Y vdd OAI21X1
XNAND3X1_5 INVX4_15/A INVX4_16/A INVX1_78/A gnd NAND3X1_6/B vdd NAND3X1
XOAI21X1_112 BUFX4_66/Y INVX1_101/A OAI21X1_112/C gnd NOR2X1_147/B vdd OAI21X1
XOAI21X1_101 INVX1_59/Y MUX2X1_27/S OAI21X1_101/C gnd OAI21X1_109/B vdd OAI21X1
XOAI21X1_167 AOI22X1_1/Y NOR2X1_120/A AOI21X1_56/Y gnd AOI21X1_57/C vdd OAI21X1
XOAI21X1_145 MUX2X1_36/A BUFX4_16/Y OAI21X1_145/C gnd MUX2X1_21/B vdd OAI21X1
XOAI21X1_134 BUFX4_35/Y MUX2X1_36/B OAI21X1_134/C gnd MUX2X1_21/A vdd OAI21X1
XOAI21X1_178 NOR2X1_83/A MUX2X1_22/Y OAI21X1_178/C gnd OAI21X1_178/Y vdd OAI21X1
XOAI21X1_156 XOR2X1_3/Y NOR2X1_112/Y AOI21X1_48/A gnd AOI21X1_51/B vdd OAI21X1
XOAI21X1_189 INVX1_89/Y BUFX4_131/Y OAI21X1_189/C gnd OAI21X1_375/B vdd OAI21X1
XINVX1_209 INVX1_209/A gnd INVX1_209/Y vdd INVX1
XOAI21X1_123 OAI21X1_123/A MUX2X1_32/S INVX8_7/A gnd AOI21X1_40/C vdd OAI21X1
XNAND2X1_173 BUFX4_46/Y operand_A[50] gnd OAI21X1_511/C vdd NAND2X1
XNAND2X1_151 operand_A[30] BUFX4_50/Y gnd OAI21X1_106/C vdd NAND2X1
XNAND2X1_184 BUFX4_191/Y OAI21X1_140/Y gnd OAI21X1_141/C vdd NAND2X1
XNAND2X1_162 BUFX4_48/Y operand_A[12] gnd OAI21X1_118/C vdd NAND2X1
XNAND2X1_195 operand_A[5] BUFX4_82/Y gnd OAI21X1_158/C vdd NAND2X1
XNAND2X1_140 MUX2X1_1/S operand_A[16] gnd OAI21X1_95/C vdd NAND2X1
XAOI22X1_18 BUFX4_58/Y AND2X2_26/B BUFX4_5/Y INVX1_202/Y gnd AOI22X1_18/Y vdd AOI22X1
XAOI22X1_29 NOR2X1_115/Y AOI22X1_29/B AOI22X1_29/C NOR2X1_59/Y gnd AOI22X1_29/Y vdd
+ AOI22X1
XOAI21X1_690 INVX4_7/Y BUFX4_46/Y OAI21X1_53/C gnd MUX2X1_76/A vdd OAI21X1
XXNOR2X1_40 XNOR2X1_40/A XOR2X1_5/Y gnd XNOR2X1_40/Y vdd XNOR2X1
XBUFX2_50 BUFX2_50/A gnd result[47] vdd BUFX2
XBUFX2_61 BUFX2_61/A gnd result[58] vdd BUFX2
XAOI21X1_73 BUFX4_148/Y INVX4_17/Y OAI22X1_3/Y gnd NAND3X1_10/B vdd AOI21X1
XAOI21X1_84 AOI21X1_84/A NOR2X1_156/Y NOR2X1_157/Y gnd AOI21X1_84/Y vdd AOI21X1
XAOI21X1_95 NAND3X1_9/A XNOR2X1_32/Y AOI21X1_95/C gnd AOI21X1_96/B vdd AOI21X1
XAOI21X1_62 AOI22X1_4/C AOI21X1_62/B BUFX4_95/Y gnd AOI21X1_64/B vdd AOI21X1
XOAI21X1_2 INVX1_4/Y NOR2X1_5/Y OAI21X1_2/C gnd NOR2X1_6/A vdd OAI21X1
XAOI21X1_40 BUFX4_163/Y AND2X2_25/A AOI21X1_40/C gnd AOI21X1_41/C vdd AOI21X1
XAOI21X1_51 AND2X2_46/B AOI21X1_51/B AOI21X1_51/C gnd AOI21X1_51/Y vdd AOI21X1
XFILL_9_0_1 gnd vdd FILL
XNOR2X1_419 operand_A[38] INVX2_67/Y gnd NOR2X1_419/Y vdd NOR2X1
XNOR2X1_408 MUX2X1_4/S operand_A[0] gnd NOR2X1_409/A vdd NOR2X1
XXOR2X1_5 operand_B[7] operand_A[7] gnd XOR2X1_5/Y vdd XOR2X1
XMUX2X1_6 operand_A[35] operand_A[34] MUX2X1_6/S gnd MUX2X1_6/Y vdd MUX2X1
XCLKBUF1_7 clk gnd CLKBUF1_7/Y vdd CLKBUF1
XBUFX4_101 DFFSR_1/Q gnd BUFX4_101/Y vdd BUFX4
XBUFX4_145 INVX8_16/Y gnd BUFX4_145/Y vdd BUFX4
XNOR2X1_238 operand_B[46] INVX2_43/Y gnd INVX1_192/A vdd NOR2X1
XNOR2X1_249 OR2X2_29/B NOR2X1_249/B gnd OR2X2_30/A vdd NOR2X1
XBUFX4_156 INVX8_14/Y gnd OAI22X1_9/A vdd BUFX4
XNOR2X1_216 operand_A[44] operand_B[44] gnd NOR2X1_217/A vdd NOR2X1
XNOR2X1_205 BUFX4_184/Y INVX1_324/A gnd NOR2X1_205/Y vdd NOR2X1
XBUFX4_167 INVX8_5/Y gnd BUFX4_167/Y vdd BUFX4
XBUFX4_189 operand_B[1] gnd NOR2X1_54/A vdd BUFX4
XBUFX4_178 operand_B[4] gnd OR2X2_43/B vdd BUFX4
XBUFX4_123 INVX8_3/Y gnd NOR2X1_19/B vdd BUFX4
XBUFX4_134 operand_B[2] gnd BUFX4_134/Y vdd BUFX4
XBUFX4_112 operand_B[5] gnd BUFX4_112/Y vdd BUFX4
XNOR2X1_227 BUFX4_183/Y MUX2X1_64/B gnd NOR2X1_227/Y vdd NOR2X1
XAOI21X1_396 BUFX4_79/Y MUX2X1_126/Y INVX8_9/Y gnd OAI22X1_34/C vdd AOI21X1
XAOI21X1_352 XNOR2X1_23/Y NOR2X1_472/B BUFX4_31/Y gnd AOI21X1_359/B vdd AOI21X1
XAOI21X1_363 NOR2X1_39/Y BUFX4_152/Y BUFX4_11/Y gnd NAND2X1_626/A vdd AOI21X1
XAOI21X1_330 NAND2X1_609/Y OAI21X1_796/Y BUFX4_112/Y gnd OAI21X1_800/B vdd AOI21X1
XAOI21X1_341 BUFX4_85/Y NOR2X1_213/Y NAND2X1_618/Y gnd NAND2X1_619/A vdd AOI21X1
XAOI21X1_385 BUFX4_78/Y OAI21X1_894/Y INVX8_9/Y gnd OAI22X1_31/B vdd AOI21X1
XINVX8_9 INVX8_9/A gnd INVX8_9/Y vdd INVX8
XAOI21X1_374 OR2X2_47/B NOR2X1_486/Y OAI21X1_874/Y gnd NOR2X1_489/A vdd AOI21X1
XDFFPOSX1_40 BUFX2_42/A CLKBUF1_3/Y DFFPOSX1_40/D gnd vdd DFFPOSX1
XDFFPOSX1_51 BUFX2_53/A CLKBUF1_4/Y DFFPOSX1_51/D gnd vdd DFFPOSX1
XDFFPOSX1_62 BUFX2_64/A CLKBUF1_5/Y DFFPOSX1_62/D gnd vdd DFFPOSX1
XBUFX4_29 INVX8_6/Y gnd BUFX4_29/Y vdd BUFX4
XBUFX4_18 INVX8_2/Y gnd BUFX4_18/Y vdd BUFX4
XFILL_22_1 gnd vdd FILL
XOAI21X1_519 INVX2_78/A INVX1_216/Y NOR2X1_280/Y gnd NAND3X1_31/C vdd OAI21X1
XOAI21X1_508 OR2X2_19/B NOR2X1_487/B OAI21X1_508/C gnd OAI21X1_508/Y vdd OAI21X1
XNAND2X1_525 INVX4_25/A OAI21X1_626/Y gnd NAND3X1_39/C vdd NAND2X1
XNAND2X1_503 BUFX4_167/Y OAI21X1_406/Y gnd NAND2X1_503/Y vdd NAND2X1
XNAND2X1_536 NOR2X1_403/Y NOR2X1_406/Y gnd NOR2X1_407/B vdd NAND2X1
XNAND2X1_514 MUX2X1_32/S OAI21X1_435/B gnd OAI21X1_605/C vdd NAND2X1
XNAND2X1_547 operand_B[36] INVX2_44/Y gnd OAI21X1_664/B vdd NAND2X1
XNAND2X1_558 BUFX4_192/Y INVX1_284/Y gnd OAI21X1_678/C vdd NAND2X1
XNAND2X1_569 BUFX4_131/Y OAI21X1_703/Y gnd OAI21X1_706/C vdd NAND2X1
XFILL_25_5_0 gnd vdd FILL
XFILL_0_5_0 gnd vdd FILL
XAOI21X1_171 INVX1_204/Y NOR2X1_259/Y BUFX4_32/Y gnd OAI21X1_488/C vdd AOI21X1
XAOI21X1_193 INVX2_78/Y OAI21X1_532/C BUFX4_93/Y gnd OAI21X1_522/C vdd AOI21X1
XAOI21X1_182 BUFX4_153/Y NOR2X1_273/A OAI22X1_9/Y gnd AND2X2_31/A vdd AOI21X1
XAOI21X1_160 NOR2X1_75/A AND2X2_7/Y NOR2X1_239/Y gnd NOR2X1_478/B vdd AOI21X1
XFILL_16_5_0 gnd vdd FILL
XOAI21X1_305 OAI21X1_305/A AOI21X1_83/Y BUFX4_101/Y gnd OAI21X1_306/C vdd OAI21X1
XOAI21X1_327 INVX2_65/A INVX2_63/A OAI21X1_327/C gnd INVX1_142/A vdd OAI21X1
XOAI21X1_316 BUFX4_61/Y OAI21X1_327/C AOI22X1_8/Y gnd NOR2X1_167/B vdd OAI21X1
XOAI21X1_349 INVX1_140/Y BUFX4_68/Y OAI21X1_349/C gnd OAI21X1_349/Y vdd OAI21X1
XOAI21X1_338 INVX1_115/Y BUFX4_120/Y OAI21X1_338/C gnd INVX1_187/A vdd OAI21X1
XBUFX4_3 BUFX4_6/A gnd BUFX4_3/Y vdd BUFX4
XNAND2X1_355 NOR2X1_174/A NAND2X1_355/B gnd INVX1_148/A vdd NAND2X1
XNAND2X1_344 INVX4_19/A INVX2_65/Y gnd OAI21X1_328/B vdd NAND2X1
XNAND2X1_322 OAI21X1_289/Y NOR2X1_162/Y gnd OAI21X1_305/A vdd NAND2X1
XNAND2X1_377 BUFX4_53/Y operand_A[40] gnd OAI21X1_382/C vdd NAND2X1
XNAND2X1_311 MUX2X1_9/S operand_A[35] gnd OAI21X1_293/C vdd NAND2X1
XNAND2X1_366 BUFX4_25/Y INVX1_88/Y gnd OAI21X1_365/C vdd NAND2X1
XNAND2X1_333 BUFX4_38/Y MUX2X1_35/Y gnd OAI21X1_320/C vdd NAND2X1
XNAND2X1_300 BUFX4_19/Y OAI21X1_415/B gnd OAI21X1_278/C vdd NAND2X1
XNAND2X1_399 AND2X2_17/B NOR2X1_218/Y gnd NOR2X1_247/B vdd NAND2X1
XNAND2X1_388 BUFX4_16/Y OAI21X1_247/A gnd OAI21X1_405/C vdd NAND2X1
XINVX4_3 operand_A[22] gnd INVX4_3/Y vdd INVX4
XOAI21X1_850 AND2X2_62/Y AND2X2_64/Y INVX8_10/A gnd NAND3X1_66/C vdd OAI21X1
XOAI21X1_861 NOR2X1_477/Y OAI21X1_862/B BUFX4_91/Y gnd NAND3X1_69/B vdd OAI21X1
XOAI21X1_883 operand_B[19] operand_A[19] BUFX4_1/Y gnd OAI21X1_884/C vdd OAI21X1
XOAI21X1_894 BUFX4_164/Y MUX2X1_34/B OAI21X1_894/C gnd OAI21X1_894/Y vdd OAI21X1
XOAI21X1_872 OAI21X1_872/A OAI21X1_872/B AND2X2_70/Y gnd OAI21X1_872/Y vdd OAI21X1
XFILL_31_3_0 gnd vdd FILL
XNAND3X1_6 INVX8_6/A NAND3X1_6/B NAND3X1_6/C gnd NAND3X1_6/Y vdd NAND3X1
XOAI21X1_135 INVX2_54/Y BUFX4_53/Y OAI21X1_412/C gnd OAI21X1_135/Y vdd OAI21X1
XFILL_22_3_0 gnd vdd FILL
XOAI21X1_102 INVX4_8/Y MUX2X1_9/S OAI21X1_102/C gnd INVX1_61/A vdd OAI21X1
XOAI21X1_124 INVX4_12/Y BUFX4_53/Y OAI21X1_628/A gnd OAI21X1_125/B vdd OAI21X1
XOAI21X1_146 BUFX4_8/Y INVX1_72/Y BUFX4_99/Y gnd OR2X2_8/B vdd OAI21X1
XOAI21X1_113 INVX2_14/Y MUX2X1_4/S OAI21X1_113/C gnd OAI21X1_113/Y vdd OAI21X1
XOAI21X1_168 NOR2X1_485/B OAI21X1_168/B AOI21X1_57/Y gnd OAI21X1_169/C vdd OAI21X1
XOAI21X1_179 OAI21X1_365/B BUFX4_37/Y OAI21X1_179/C gnd INVX1_86/A vdd OAI21X1
XOAI21X1_157 XOR2X1_4/Y OAI21X1_743/C INVX1_80/Y gnd AOI21X1_51/C vdd OAI21X1
XNAND2X1_185 MUX2X1_5/S operand_A[34] gnd OAI21X1_275/C vdd NAND2X1
XNAND2X1_130 NOR2X1_54/A OAI21X1_77/Y gnd OAI21X1_78/C vdd NAND2X1
XNAND2X1_174 MUX2X1_97/S OAI21X1_129/Y gnd OAI21X1_130/C vdd NAND2X1
XNAND2X1_152 BUFX4_68/Y OAI21X1_106/Y gnd OAI21X1_107/C vdd NAND2X1
XNAND2X1_163 BUFX4_50/Y operand_A[14] gnd OAI21X1_119/C vdd NAND2X1
XNAND2X1_196 OAI21X1_158/C NAND2X1_73/Y gnd NAND3X1_4/A vdd NAND2X1
XFILL_5_4_0 gnd vdd FILL
XNAND2X1_141 MUX2X1_6/S operand_A[18] gnd OAI21X1_96/C vdd NAND2X1
XFILL_13_3_0 gnd vdd FILL
XAOI22X1_19 BUFX4_91/Y AOI22X1_19/B MUX2X1_44/Y INVX8_7/A gnd AOI22X1_19/Y vdd AOI22X1
XOAI21X1_691 INVX2_12/Y BUFX4_48/Y OAI21X1_52/C gnd NOR2X1_432/B vdd OAI21X1
XOAI21X1_680 INVX4_5/Y MUX2X1_6/S OAI21X1_39/C gnd OAI21X1_680/Y vdd OAI21X1
XXNOR2X1_30 XNOR2X1_30/A INVX4_16/Y gnd XNOR2X1_30/Y vdd XNOR2X1
XXNOR2X1_41 XNOR2X1_41/A XNOR2X1_41/B gnd XNOR2X1_41/Y vdd XNOR2X1
XBUFX2_40 BUFX2_40/A gnd result[37] vdd BUFX2
XBUFX2_51 BUFX2_51/A gnd result[48] vdd BUFX2
XBUFX2_62 BUFX2_62/A gnd result[59] vdd BUFX2
XAOI21X1_41 INVX8_9/A MUX2X1_21/Y AOI21X1_41/C gnd AOI21X1_41/Y vdd AOI21X1
XAOI21X1_30 INVX1_85/A INVX2_18/Y INVX1_30/Y gnd OAI21X1_31/C vdd AOI21X1
XAOI21X1_52 AOI21X1_52/A NOR2X1_114/Y AOI21X1_52/C gnd AOI21X1_52/Y vdd AOI21X1
XAOI21X1_96 AOI21X1_96/A AOI21X1_96/B NOR2X1_163/Y gnd AOI21X1_96/Y vdd AOI21X1
XAOI21X1_85 INVX4_19/Y INVX1_144/A BUFX4_95/Y gnd AOI21X1_85/Y vdd AOI21X1
XAOI21X1_63 INVX4_18/A INVX1_100/Y OR2X2_4/Y gnd AOI21X1_63/Y vdd AOI21X1
XAOI21X1_74 INVX8_15/A AOI21X1_74/B NAND3X1_10/Y gnd AOI21X1_74/Y vdd AOI21X1
XOAI21X1_3 OAI21X1_3/A OAI21X1_3/B OAI21X1_3/C gnd OAI21X1_3/Y vdd OAI21X1
XNOR2X1_409 NOR2X1_409/A INVX2_10/Y gnd NOR2X1_410/B vdd NOR2X1
XFILL_27_2_0 gnd vdd FILL
XFILL_2_2_0 gnd vdd FILL
XXOR2X1_6 operand_A[11] operand_B[11] gnd XOR2X1_6/Y vdd XOR2X1
XMUX2X1_7 operand_A[31] operand_A[30] MUX2X1_7/S gnd MUX2X1_7/Y vdd MUX2X1
XCLKBUF1_8 clk gnd CLKBUF1_8/Y vdd CLKBUF1
XFILL_10_1_0 gnd vdd FILL
XBUFX4_102 DFFSR_1/Q gnd BUFX4_102/Y vdd BUFX4
XBUFX4_146 INVX8_16/Y gnd OAI22X1_9/C vdd BUFX4
XBUFX4_157 INVX8_14/Y gnd BUFX4_157/Y vdd BUFX4
XNOR2X1_217 NOR2X1_217/A AND2X2_21/Y gnd INVX2_75/A vdd NOR2X1
XFILL_18_2_0 gnd vdd FILL
XNOR2X1_239 OR2X2_7/B MUX2X1_21/A gnd NOR2X1_239/Y vdd NOR2X1
XNOR2X1_206 BUFX4_36/Y INVX1_109/Y gnd NOR2X1_206/Y vdd NOR2X1
XBUFX4_124 INVX8_3/Y gnd MUX2X1_71/S vdd BUFX4
XNOR2X1_228 OR2X2_13/B NOR2X1_228/B gnd NOR2X1_228/Y vdd NOR2X1
XBUFX4_135 operand_B[2] gnd MUX2X1_87/S vdd BUFX4
XBUFX4_179 operand_B[4] gnd BUFX4_179/Y vdd BUFX4
XBUFX4_113 operand_B[5] gnd BUFX4_113/Y vdd BUFX4
XBUFX4_168 INVX8_5/Y gnd MUX2X1_25/S vdd BUFX4
XDFFPOSX1_30 BUFX2_32/A CLKBUF1_1/Y DFFPOSX1_30/D gnd vdd DFFPOSX1
XDFFPOSX1_41 BUFX2_43/A CLKBUF1_3/Y OAI21X1_378/Y gnd vdd DFFPOSX1
XDFFPOSX1_52 BUFX2_54/A CLKBUF1_4/Y DFFPOSX1_52/D gnd vdd DFFPOSX1
XDFFPOSX1_63 BUFX2_65/A CLKBUF1_5/Y DFFPOSX1_63/D gnd vdd DFFPOSX1
XAOI21X1_397 NOR2X1_42/Y BUFX4_148/Y BUFX4_13/Y gnd NAND3X1_72/B vdd AOI21X1
XAOI21X1_386 BUFX4_108/Y XNOR2X1_45/Y NAND2X1_638/Y gnd OAI21X1_898/C vdd AOI21X1
XAOI21X1_353 INVX1_82/Y INVX1_314/Y INVX1_84/Y gnd OR2X2_45/A vdd AOI21X1
XAOI21X1_331 INVX2_17/Y OAI21X1_805/B BUFX4_27/Y gnd OAI21X1_805/C vdd AOI21X1
XAOI21X1_320 INVX8_10/A OAI21X1_765/Y NOR2X1_444/Y gnd NAND3X1_62/C vdd AOI21X1
XAOI21X1_342 BUFX4_89/Y OAI21X1_829/Y NAND2X1_619/Y gnd AND2X2_60/A vdd AOI21X1
XAOI21X1_375 BUFX4_78/Y MUX2X1_124/Y INVX8_9/Y gnd OAI22X1_29/C vdd AOI21X1
XAOI21X1_364 INVX8_15/A INVX1_193/Y NAND2X1_626/Y gnd NAND3X1_69/A vdd AOI21X1
XBUFX4_19 INVX8_2/Y gnd BUFX4_19/Y vdd BUFX4
XOAI21X1_509 INVX1_212/Y NOR2X1_273/Y OAI21X1_509/C gnd OAI21X1_509/Y vdd OAI21X1
XNAND2X1_548 operand_B[34] INVX2_60/Y gnd OAI21X1_665/B vdd NAND2X1
XNAND2X1_537 INVX1_233/A NOR2X1_411/Y gnd NOR2X1_412/B vdd NAND2X1
XNAND2X1_526 operand_A[62] INVX1_256/Y gnd NAND3X1_40/B vdd NAND2X1
XINVX1_190 operand_A[47] gnd INVX1_190/Y vdd INVX1
XNAND2X1_504 MUX2X1_66/S MUX2X1_66/B gnd AOI22X1_26/A vdd NAND2X1
XNAND2X1_515 BUFX4_167/Y INVX1_176/A gnd OAI21X1_939/A vdd NAND2X1
XNAND2X1_559 MUX2X1_98/S OAI21X1_680/Y gnd OAI21X1_681/C vdd NAND2X1
XFILL_25_5_1 gnd vdd FILL
XFILL_0_5_1 gnd vdd FILL
XFILL_24_0_0 gnd vdd FILL
XAOI21X1_150 NAND3X1_9/A XNOR2X1_34/Y NAND3X1_24/Y gnd AOI21X1_151/B vdd AOI21X1
XAOI21X1_194 INVX4_20/A OAI21X1_523/Y INVX1_145/A gnd NAND2X1_469/A vdd AOI21X1
XAOI21X1_161 INVX4_18/A INVX1_193/Y NAND3X1_28/Y gnd OAI21X1_465/C vdd AOI21X1
XAOI21X1_183 BUFX4_112/Y OAI22X1_29/D OR2X2_31/Y gnd OAI21X1_508/C vdd AOI21X1
XAOI21X1_172 INVX8_4/A OAI21X1_494/Y OAI21X1_496/Y gnd OAI21X1_497/C vdd AOI21X1
XFILL_7_1_0 gnd vdd FILL
XFILL_16_5_1 gnd vdd FILL
XFILL_15_0_0 gnd vdd FILL
XOAI21X1_306 NOR2X1_93/A INVX1_125/Y OAI21X1_306/C gnd OAI21X1_306/Y vdd OAI21X1
XOAI21X1_328 INVX2_64/Y OAI21X1_328/B INVX1_142/Y gnd AOI21X1_97/B vdd OAI21X1
XOAI21X1_317 NOR2X1_444/B OR2X2_32/B NOR2X1_167/Y gnd AOI21X1_93/C vdd OAI21X1
XBUFX4_4 BUFX4_6/A gnd BUFX4_4/Y vdd BUFX4
XOAI21X1_339 INVX1_42/Y BUFX4_17/Y OAI21X1_339/C gnd OAI21X1_339/Y vdd OAI21X1
XNAND2X1_356 INVX2_68/Y AOI21X1_97/B gnd OAI21X1_346/C vdd NAND2X1
XNAND2X1_345 OAI21X1_329/Y AOI22X1_9/Y gnd OAI21X1_344/A vdd NAND2X1
XNAND2X1_323 operand_A[37] operand_B[37] gnd OAI21X1_327/C vdd NAND2X1
XNAND2X1_389 INVX1_169/A OAI21X1_393/B gnd OAI21X1_408/C vdd NAND2X1
XNAND2X1_378 NOR2X1_54/A OAI21X1_348/Y gnd OAI21X1_383/C vdd NAND2X1
XNAND2X1_312 MUX2X1_97/S OAI21X1_257/Y gnd OAI21X1_294/C vdd NAND2X1
XNAND2X1_367 BUFX4_163/Y MUX2X1_126/A gnd OAI21X1_366/C vdd NAND2X1
XNAND2X1_301 MUX2X1_49/S MUX2X1_46/B gnd OAI21X1_282/C vdd NAND2X1
XNAND2X1_334 BUFX4_122/Y OAI21X1_219/Y gnd OAI21X1_321/C vdd NAND2X1
XOAI21X1_862 NOR2X1_478/Y OAI21X1_862/B INVX8_10/A gnd NAND3X1_69/C vdd OAI21X1
XINVX4_4 operand_A[21] gnd INVX4_4/Y vdd INVX4
XOAI21X1_851 INVX2_18/Y INVX2_19/Y OR2X2_45/A gnd NAND3X1_67/B vdd OAI21X1
XOAI21X1_840 INVX8_15/Y INVX1_310/Y OAI21X1_840/C gnd NOR2X1_468/B vdd OAI21X1
XOAI21X1_884 BUFX4_65/Y INVX1_319/Y OAI21X1_884/C gnd NOR2X1_490/B vdd OAI21X1
XOAI21X1_873 INVX1_315/Y OAI21X1_7/Y OAI21X1_3/B gnd OR2X2_47/A vdd OAI21X1
XOAI21X1_895 operand_B[21] operand_A[21] BUFX4_3/Y gnd OAI21X1_896/C vdd OAI21X1
XFILL_31_3_1 gnd vdd FILL
XNAND3X1_7 NOR2X1_19/B OR2X2_39/B NAND3X1_7/C gnd NAND3X1_7/Y vdd NAND3X1
XOAI21X1_147 BUFX4_158/Y OAI21X1_94/C AOI22X1_3/Y gnd AOI21X1_42/C vdd OAI21X1
XOAI21X1_169 INVX4_15/Y NOR2X1_103/A OAI21X1_169/C gnd AOI21X1_64/A vdd OAI21X1
XFILL_22_3_1 gnd vdd FILL
XOAI21X1_103 INVX2_30/Y MUX2X1_5/S OAI21X1_704/C gnd OAI21X1_103/Y vdd OAI21X1
XOAI21X1_136 XOR2X1_3/A MUX2X1_17/Y OAI21X1_136/C gnd INVX1_70/A vdd OAI21X1
XOAI21X1_125 BUFX4_69/Y OAI21X1_125/B OAI21X1_125/C gnd OAI21X1_272/A vdd OAI21X1
XOAI21X1_158 NOR2X1_23/Y NAND2X1_26/A OAI21X1_158/C gnd AOI21X1_52/A vdd OAI21X1
XOAI21X1_114 XOR2X1_3/A MUX2X1_11/Y OAI21X1_114/C gnd INVX1_122/A vdd OAI21X1
XBUFX2_1 gnd gnd carry_flag vdd BUFX2
XNAND2X1_197 NOR2X1_3/Y AND2X2_9/A gnd NOR2X1_110/A vdd NAND2X1
XNAND2X1_175 MUX2X1_1/S operand_A[54] gnd OAI21X1_556/C vdd NAND2X1
XNAND2X1_186 MUX2X1_1/S operand_A[32] gnd OAI21X1_217/C vdd NAND2X1
XNAND2X1_131 BUFX4_43/Y operand_A[45] gnd OAI21X1_80/C vdd NAND2X1
XNAND2X1_120 BUFX4_68/Y INVX1_48/Y gnd OAI21X1_69/C vdd NAND2X1
XNAND2X1_164 BUFX4_74/Y INVX1_102/A gnd OAI21X1_120/C vdd NAND2X1
XNAND2X1_142 BUFX4_76/Y OAI21X1_96/Y gnd OAI21X1_97/C vdd NAND2X1
XFILL_5_4_1 gnd vdd FILL
XNAND2X1_153 BUFX4_122/Y OAI21X1_107/Y gnd OAI21X1_108/C vdd NAND2X1
XINVX2_1 operand_B[29] gnd INVX2_1/Y vdd INVX2
XFILL_13_3_1 gnd vdd FILL
XAOI21X1_1 NOR2X1_2/Y NAND2X1_3/Y NOR2X1_1/Y gnd INVX1_2/A vdd AOI21X1
XOAI21X1_670 operand_A[42] INVX2_72/Y NAND3X1_21/C gnd OAI21X1_671/C vdd OAI21X1
XOAI21X1_692 NOR2X1_432/B BUFX4_66/Y NOR2X1_19/B gnd OAI21X1_692/Y vdd OAI21X1
XOAI21X1_681 INVX1_285/Y NOR2X1_82/A OAI21X1_681/C gnd MUX2X1_74/B vdd OAI21X1
XXNOR2X1_31 XNOR2X1_31/A INVX2_62/Y gnd XNOR2X1_31/Y vdd XNOR2X1
XXNOR2X1_20 BUFX4_112/Y operand_A[5] gnd XNOR2X1_20/Y vdd XNOR2X1
XXNOR2X1_42 XNOR2X1_42/A INVX4_26/Y gnd XNOR2X1_42/Y vdd XNOR2X1
XBUFX2_41 OR2X2_36/A gnd result[38] vdd BUFX2
XBUFX2_52 BUFX2_52/A gnd result[49] vdd BUFX2
XBUFX2_63 BUFX2_63/A gnd result[60] vdd BUFX2
XBUFX2_30 BUFX2_30/A gnd result[27] vdd BUFX2
XAOI21X1_64 AOI21X1_64/A AOI21X1_64/B OR2X2_5/Y gnd AOI21X1_65/B vdd AOI21X1
XAOI21X1_42 OR2X2_40/B INVX1_74/Y AOI21X1_42/C gnd AND2X2_8/A vdd AOI21X1
XAOI21X1_86 XOR2X1_4/A INVX1_118/A INVX1_133/A gnd AOI21X1_86/Y vdd AOI21X1
XAOI21X1_20 INVX1_4/A NOR2X1_52/Y NOR2X1_5/Y gnd OAI21X1_27/B vdd AOI21X1
XAOI21X1_75 BUFX4_83/Y AOI21X1_75/B AOI21X1_75/C gnd AND2X2_13/A vdd AOI21X1
XAOI21X1_31 NOR2X1_59/Y OAI21X1_30/Y OAI21X1_31/Y gnd OAI21X1_32/C vdd AOI21X1
XAOI21X1_53 AOI21X1_53/A NOR2X1_116/Y AOI21X1_53/C gnd AOI21X1_53/Y vdd AOI21X1
XAOI21X1_97 INVX2_68/Y AOI21X1_97/B BUFX4_28/Y gnd AOI21X1_97/Y vdd AOI21X1
XOAI21X1_4 INVX2_3/Y INVX2_4/Y OAI21X1_4/C gnd OAI21X1_5/C vdd OAI21X1
XFILL_3_1 gnd vdd FILL
XFILL_27_2_1 gnd vdd FILL
XFILL_2_2_1 gnd vdd FILL
XXOR2X1_7 XOR2X1_7/A operand_A[2] gnd XOR2X1_7/Y vdd XOR2X1
XMUX2X1_8 operand_A[43] operand_A[42] MUX2X1_8/S gnd MUX2X1_8/Y vdd MUX2X1
XFILL_10_1_1 gnd vdd FILL
XBUFX4_103 DFFSR_1/Q gnd NOR2X1_93/A vdd BUFX4
XBUFX4_136 operand_B[2] gnd BUFX4_136/Y vdd BUFX4
XBUFX4_125 INVX8_3/Y gnd BUFX4_125/Y vdd BUFX4
XBUFX4_114 operand_B[5] gnd BUFX4_114/Y vdd BUFX4
XNOR2X1_207 BUFX4_101/Y BUFX2_45/A gnd NOR2X1_207/Y vdd NOR2X1
XBUFX4_147 INVX8_16/Y gnd OAI22X1_3/C vdd BUFX4
XNOR2X1_218 INVX1_169/A INVX2_74/A gnd NOR2X1_218/Y vdd NOR2X1
XBUFX4_158 INVX8_14/Y gnd BUFX4_158/Y vdd BUFX4
XNOR2X1_229 INVX2_43/Y INVX1_184/Y gnd NOR2X1_231/B vdd NOR2X1
XFILL_18_2_1 gnd vdd FILL
XBUFX4_169 INVX8_10/Y gnd BUFX4_169/Y vdd BUFX4
XAOI21X1_343 NOR2X1_60/Y AOI21X1_55/B OAI21X1_30/Y gnd INVX1_314/A vdd AOI21X1
XAOI21X1_321 BUFX4_82/Y OAI22X1_6/B OR2X2_41/Y gnd OAI21X1_777/C vdd AOI21X1
XAOI21X1_332 INVX2_17/A OAI21X1_807/A OAI21X1_807/Y gnd NOR2X1_454/A vdd AOI21X1
XAOI21X1_310 NOR2X1_75/A INVX1_318/A OAI21X1_740/Y gnd NOR2X1_438/A vdd AOI21X1
XDFFPOSX1_53 BUFX2_55/A CLKBUF1_4/Y OAI21X1_530/Y gnd vdd DFFPOSX1
XDFFPOSX1_31 BUFX2_33/A CLKBUF1_1/Y AOI21X1_37/Y gnd vdd DFFPOSX1
XDFFPOSX1_42 OR2X2_36/B CLKBUF1_8/Y DFFPOSX1_42/D gnd vdd DFFPOSX1
XDFFPOSX1_64 BUFX2_66/A CLKBUF1_5/Y DFFPOSX1_64/D gnd vdd DFFPOSX1
XAOI21X1_398 OAI21X1_909/Y NOR2X1_499/Y NOR2X1_498/Y gnd DFFPOSX1_25/D vdd AOI21X1
XAOI21X1_387 INVX2_94/A OAI21X1_902/B BUFX4_96/Y gnd OAI21X1_902/C vdd AOI21X1
XAOI21X1_354 BUFX4_41/Y MUX2X1_112/A BUFX4_183/Y gnd OAI21X1_852/C vdd AOI21X1
XAOI21X1_365 NOR2X1_479/Y OAI21X1_857/Y NOR2X1_480/Y gnd DFFPOSX1_16/D vdd AOI21X1
XAOI21X1_376 XOR2X1_2/Y OAI21X1_880/B BUFX4_31/Y gnd OAI21X1_880/C vdd AOI21X1
XDFFPOSX1_20 BUFX2_22/A DFFSR_1/CLK AOI22X1_49/Y gnd vdd DFFPOSX1
XNAND2X1_516 OAI21X1_622/C BUFX4_143/Y gnd NAND2X1_516/Y vdd NAND2X1
XNAND2X1_549 operand_B[33] INVX2_56/Y gnd OAI21X1_666/C vdd NAND2X1
XINVX1_191 operand_B[47] gnd INVX1_191/Y vdd INVX1
XNAND2X1_527 operand_A[63] INVX8_12/A gnd NAND3X1_41/A vdd NAND2X1
XINVX1_180 INVX1_180/A gnd INVX1_180/Y vdd INVX1
XNAND2X1_538 NOR2X1_122/Y NOR2X1_412/Y gnd NOR2X1_413/B vdd NAND2X1
XNAND2X1_505 BUFX4_167/Y NOR2X1_206/Y gnd OAI21X1_926/A vdd NAND2X1
XFILL_24_0_1 gnd vdd FILL
XAOI21X1_184 INVX8_11/A XNOR2X1_37/Y OAI21X1_508/Y gnd AOI21X1_185/B vdd AOI21X1
XAOI21X1_173 INVX8_11/A XNOR2X1_36/Y OAI21X1_497/Y gnd AOI21X1_174/A vdd AOI21X1
XAOI21X1_140 NOR2X1_202/B INVX2_74/A NOR2X1_210/B gnd OAI21X1_424/C vdd AOI21X1
XAOI21X1_162 BUFX4_107/Y XNOR2X1_35/Y OR2X2_27/Y gnd AOI21X1_163/A vdd AOI21X1
XAOI21X1_151 OAI21X1_437/Y AOI21X1_151/B NOR2X1_225/Y gnd DFFPOSX1_46/D vdd AOI21X1
XAOI21X1_195 INVX1_219/Y NOR2X1_286/Y BUFX4_32/Y gnd OAI21X1_531/C vdd AOI21X1
XFILL_7_1_1 gnd vdd FILL
XFILL_15_0_1 gnd vdd FILL
XOAI21X1_329 INVX2_68/Y AOI21X1_97/B AOI21X1_97/Y gnd OAI21X1_329/Y vdd OAI21X1
XOAI21X1_307 INVX2_65/A AOI21X1_90/B AOI21X1_90/Y gnd AOI21X1_96/A vdd OAI21X1
XOAI21X1_318 BUFX4_22/Y NOR2X1_228/B INVX1_135/Y gnd MUX2X1_34/A vdd OAI21X1
XBUFX4_5 BUFX4_6/A gnd BUFX4_5/Y vdd BUFX4
XNAND2X1_302 MUX2X1_2/S INVX1_67/A gnd OAI21X1_279/C vdd NAND2X1
XNAND2X1_324 OAI21X1_327/C OR2X2_11/Y gnd INVX2_65/A vdd NAND2X1
XNAND2X1_368 MUX2X1_6/S operand_A[39] gnd OAI21X1_371/C vdd NAND2X1
XNAND2X1_335 MUX2X1_5/S operand_A[36] gnd OAI21X1_322/C vdd NAND2X1
XNAND2X1_357 BUFX4_68/Y OAI21X1_348/Y gnd OAI21X1_349/C vdd NAND2X1
XNAND2X1_379 INVX8_3/A OAI21X1_323/Y gnd OAI21X1_384/C vdd NAND2X1
XNAND2X1_313 BUFX4_136/Y OAI21X1_199/Y gnd OAI21X1_295/C vdd NAND2X1
XNAND2X1_346 BUFX4_25/Y OAI21X1_84/Y gnd OAI21X1_332/C vdd NAND2X1
XNOR2X1_390 BUFX2_58/A BUFX2_59/A gnd NOR2X1_390/Y vdd NOR2X1
XOAI21X1_896 BUFX4_155/Y AND2X2_71/B OAI21X1_896/C gnd NOR2X1_495/B vdd OAI21X1
XOAI21X1_830 AND2X2_59/Y NOR2X1_462/Y INVX8_10/A gnd OAI21X1_830/Y vdd OAI21X1
XINVX4_5 operand_A[18] gnd INVX4_5/Y vdd INVX4
XOAI21X1_863 OAI21X1_7/C INVX1_315/A NOR2X1_482/Y gnd AND2X2_67/A vdd OAI21X1
XOAI21X1_852 BUFX4_42/Y OAI21X1_852/B OAI21X1_852/C gnd OAI21X1_852/Y vdd OAI21X1
XOAI21X1_841 BUFX4_7/Y OAI21X1_841/B NOR2X1_468/Y gnd OAI21X1_842/A vdd OAI21X1
XOAI21X1_885 BUFX4_155/Y XNOR2X1_15/Y BUFX4_100/Y gnd NOR2X1_490/A vdd OAI21X1
XOAI21X1_874 NOR2X1_486/Y OR2X2_47/B BUFX4_138/Y gnd OAI21X1_874/Y vdd OAI21X1
XNAND3X1_8 NAND3X1_8/A NAND3X1_8/B NAND3X1_8/C gnd NAND3X1_8/Y vdd NAND3X1
XOAI21X1_126 INVX4_13/Y MUX2X1_4/S OAI21X1_591/C gnd OAI21X1_126/Y vdd OAI21X1
XOAI21X1_137 INVX4_14/Y BUFX4_43/Y OAI21X1_467/C gnd OAI21X1_223/B vdd OAI21X1
XOAI21X1_148 AOI21X1_41/Y BUFX4_116/Y AND2X2_8/Y gnd AOI21X1_43/C vdd OAI21X1
XOAI21X1_159 NOR2X1_21/Y NAND2X1_23/A INVX1_81/Y gnd AOI21X1_52/C vdd OAI21X1
XOAI21X1_115 NOR2X1_147/B BUFX4_125/Y OAI21X1_115/C gnd INVX1_66/A vdd OAI21X1
XOAI21X1_104 INVX1_61/Y BUFX4_67/Y OAI21X1_104/C gnd INVX1_62/A vdd OAI21X1
XNAND2X1_121 MUX2X1_9/S operand_A[49] gnd OAI21X1_70/C vdd NAND2X1
XNAND2X1_132 BUFX4_191/Y OAI21X1_80/Y gnd OAI21X1_81/C vdd NAND2X1
XBUFX2_2 gnd gnd overflow_flag vdd BUFX2
XNAND2X1_143 BUFX4_53/Y operand_A[20] gnd OAI21X1_98/C vdd NAND2X1
XNAND2X1_110 BUFX4_183/Y INVX8_7/A gnd OAI22X1_1/B vdd NAND2X1
XNAND2X1_187 BUFX4_72/Y OAI21X1_703/B gnd OAI21X1_144/C vdd NAND2X1
XNAND2X1_198 AND2X2_1/Y NOR2X1_110/Y gnd AOI21X1_50/C vdd NAND2X1
XNAND2X1_176 NOR2X1_82/A OAI21X1_229/B gnd OAI21X1_132/C vdd NAND2X1
XNAND2X1_165 MUX2X1_2/S OAI21X1_120/Y gnd OAI21X1_121/C vdd NAND2X1
XNAND2X1_154 BUFX4_23/Y INVX1_64/Y gnd OAI21X1_109/C vdd NAND2X1
XINVX2_2 operand_A[29] gnd INVX2_2/Y vdd INVX2
XOAI21X1_660 INVX2_79/A OAI21X1_660/B OAI21X1_660/C gnd OAI21X1_660/Y vdd OAI21X1
XOAI21X1_671 INVX2_73/Y operand_B[43] OAI21X1_671/C gnd OAI21X1_671/Y vdd OAI21X1
XOAI21X1_682 INVX2_26/Y BUFX4_53/Y OAI21X1_682/C gnd INVX1_286/A vdd OAI21X1
XOAI21X1_693 NOR2X1_425/Y OAI21X1_693/B OR2X2_39/B gnd NAND3X1_56/B vdd OAI21X1
XAOI21X1_2 AOI21X1_2/A OR2X2_46/B NOR2X1_7/Y gnd OAI21X1_3/B vdd AOI21X1
XXNOR2X1_32 XNOR2X1_32/A INVX2_65/A gnd XNOR2X1_32/Y vdd XNOR2X1
XXNOR2X1_10 operand_B[22] operand_A[22] gnd INVX2_94/A vdd XNOR2X1
XXNOR2X1_21 MUX2X1_34/S operand_A[4] gnd XNOR2X1_21/Y vdd XNOR2X1
XXNOR2X1_43 XNOR2X1_43/A XOR2X1_2/Y gnd XNOR2X1_43/Y vdd XNOR2X1
XBUFX2_42 BUFX2_42/A gnd result[39] vdd BUFX2
XBUFX2_53 BUFX2_53/A gnd result[50] vdd BUFX2
XBUFX2_64 BUFX2_64/A gnd result[61] vdd BUFX2
XBUFX2_31 BUFX2_31/A gnd result[28] vdd BUFX2
XBUFX2_20 BUFX2_20/A gnd result[17] vdd BUFX2
XAOI21X1_76 AOI21X1_76/A AND2X2_13/Y NOR2X1_143/Y gnd AOI21X1_76/Y vdd AOI21X1
XAOI21X1_43 OAI21X1_94/Y AOI21X1_43/B AOI21X1_43/C gnd AOI21X1_44/A vdd AOI21X1
XAOI21X1_98 NOR2X1_164/Y INVX2_65/A NOR2X1_169/Y gnd NOR2X1_183/A vdd AOI21X1
XAOI21X1_65 AOI21X1_65/A AOI21X1_65/B NOR2X1_130/Y gnd AOI21X1_65/Y vdd AOI21X1
XAOI21X1_87 INVX4_20/A AND2X2_55/A INVX1_145/A gnd NAND3X1_12/C vdd AOI21X1
XAOI21X1_32 INVX1_31/Y OAI21X1_32/Y NAND2X1_66/Y gnd OAI21X1_34/A vdd AOI21X1
XAOI21X1_21 NAND2X1_65/Y NOR2X1_4/Y NOR2X1_53/Y gnd OAI21X1_27/C vdd AOI21X1
XOAI21X1_5 operand_B[21] operand_A[21] OAI21X1_5/C gnd OAI21X1_6/B vdd OAI21X1
XAOI21X1_54 NOR2X1_115/Y INVX1_84/Y AOI21X1_54/C gnd AOI21X1_54/Y vdd AOI21X1
XAOI21X1_10 NAND2X1_41/Y NOR2X1_33/Y NOR2X1_32/Y gnd OAI21X1_17/B vdd AOI21X1
XOAI21X1_490 MUX2X1_29/Y OR2X2_43/B INVX4_11/Y gnd AOI22X1_19/B vdd OAI21X1
XFILL_3_2 gnd vdd FILL
XXOR2X1_8 operand_B[10] operand_A[10] gnd XOR2X1_8/Y vdd XOR2X1
XMUX2X1_9 operand_A[39] operand_A[38] MUX2X1_9/S gnd MUX2X1_9/Y vdd MUX2X1
XBUFX4_104 DFFSR_1/Q gnd OR2X2_48/A vdd BUFX4
XBUFX4_148 NOR2X1_89/Y gnd BUFX4_148/Y vdd BUFX4
XBUFX4_126 INVX8_3/Y gnd MUX2X1_62/S vdd BUFX4
XBUFX4_159 INVX8_5/Y gnd BUFX4_159/Y vdd BUFX4
XBUFX4_137 operand_B[2] gnd XOR2X1_7/A vdd BUFX4
XBUFX4_115 operand_B[5] gnd OR2X2_40/B vdd BUFX4
XNOR2X1_219 NOR2X1_219/A NOR2X1_219/B gnd NOR2X1_219/Y vdd NOR2X1
XNOR2X1_208 operand_A[43] operand_B[43] gnd OAI22X1_7/D vdd NOR2X1
XFILL_20_4_0 gnd vdd FILL
XAOI21X1_344 NAND2X1_40/B INVX1_314/A OAI21X1_834/Y gnd AOI21X1_345/C vdd AOI21X1
XAOI21X1_311 XOR2X1_4/Y OAI21X1_742/B BUFX4_27/Y gnd OAI21X1_742/C vdd AOI21X1
XAOI21X1_333 NAND2X1_41/Y BUFX4_1/Y BUFX4_14/Y gnd NAND3X1_63/A vdd AOI21X1
XAOI21X1_322 BUFX4_90/Y OAI21X1_771/Y OAI21X1_777/Y gnd AOI21X1_325/A vdd AOI21X1
XAOI21X1_300 INVX8_9/A OAI21X1_695/Y OAI21X1_698/Y gnd AOI22X1_31/D vdd AOI21X1
XAOI21X1_366 OAI21X1_7/C NOR2X1_485/B OAI21X1_864/Y gnd NOR2X1_483/B vdd AOI21X1
XAOI21X1_355 OAI21X1_852/Y NAND2X1_623/Y BUFX4_113/Y gnd OAI21X1_853/B vdd AOI21X1
XDFFPOSX1_54 BUFX2_56/A CLKBUF1_4/Y DFFPOSX1_54/D gnd vdd DFFPOSX1
XDFFPOSX1_32 BUFX2_34/A CLKBUF1_3/Y AOI21X1_44/Y gnd vdd DFFPOSX1
XDFFPOSX1_43 BUFX2_45/A CLKBUF1_8/Y DFFPOSX1_43/D gnd vdd DFFPOSX1
XAOI21X1_399 NAND2X1_59/A OAI21X1_915/A OAI21X1_915/Y gnd OAI21X1_919/B vdd AOI21X1
XAOI21X1_388 BUFX4_79/Y MUX2X1_125/Y INVX8_9/Y gnd OAI22X1_32/C vdd AOI21X1
XDFFPOSX1_21 BUFX2_23/A DFFSR_1/CLK OAI21X1_890/Y gnd vdd DFFPOSX1
XDFFPOSX1_10 BUFX2_12/A CLKBUF1_2/Y AOI22X1_39/Y gnd vdd DFFPOSX1
XAOI21X1_377 BUFX4_78/Y OAI21X1_882/Y INVX8_9/Y gnd OAI22X1_30/C vdd AOI21X1
XFILL_28_5_0 gnd vdd FILL
XFILL_3_5_0 gnd vdd FILL
XFILL_11_4_0 gnd vdd FILL
XFILL_19_5_0 gnd vdd FILL
XINVX1_170 INVX1_170/A gnd INVX1_170/Y vdd INVX1
XNAND2X1_506 OR2X2_34/B NOR2X1_341/Y gnd NAND3X1_35/C vdd NAND2X1
XNAND2X1_528 AND2X2_44/Y BUFX4_149/Y gnd OAI21X1_635/C vdd NAND2X1
XINVX1_192 INVX1_192/A gnd INVX1_192/Y vdd INVX1
XNAND2X1_517 BUFX4_53/Y operand_A[60] gnd OAI21X1_613/C vdd NAND2X1
XINVX1_181 INVX1_181/A gnd INVX1_181/Y vdd INVX1
XNAND2X1_539 operand_B[8] INVX2_26/Y gnd INVX1_278/A vdd NAND2X1
XAOI21X1_185 OAI21X1_498/Y AOI21X1_185/B NOR2X1_260/Y gnd DFFPOSX1_51/D vdd AOI21X1
XAOI21X1_174 AOI21X1_174/A OAI21X1_488/Y NOR2X1_255/Y gnd DFFPOSX1_50/D vdd AOI21X1
XAOI21X1_130 NAND2X1_384/Y AND2X2_19/Y NAND3X1_19/Y gnd AOI21X1_131/B vdd AOI21X1
XAOI21X1_163 AOI21X1_163/A NAND3X1_27/Y NOR2X1_237/Y gnd DFFPOSX1_48/D vdd AOI21X1
XAOI21X1_152 INVX1_186/A OAI21X1_453/B BUFX4_28/Y gnd OAI21X1_453/C vdd AOI21X1
XAOI21X1_141 NOR2X1_219/Y INVX1_155/A OAI21X1_424/Y gnd NOR2X1_220/B vdd AOI21X1
XAOI21X1_196 BUFX4_164/Y INVX1_221/Y INVX4_11/A gnd NOR2X1_493/B vdd AOI21X1
XFILL_20_1 gnd vdd FILL
XOAI21X1_308 BUFX4_122/Y OAI21X1_308/B OAI21X1_308/C gnd INVX1_183/A vdd OAI21X1
XOAI21X1_319 INVX1_136/Y MUX2X1_27/S OAI21X1_319/C gnd INVX1_137/A vdd OAI21X1
XBUFX4_6 BUFX4_6/A gnd BUFX4_6/Y vdd BUFX4
XNAND2X1_336 INVX8_1/A OAI21X1_275/Y gnd OAI21X1_323/C vdd NAND2X1
XNAND2X1_325 BUFX4_122/Y OAI21X1_225/B gnd OAI21X1_308/C vdd NAND2X1
XNAND2X1_314 BUFX4_18/Y MUX2X1_40/B gnd OAI21X1_296/C vdd NAND2X1
XNAND2X1_303 MUX2X1_51/S OAI21X1_120/Y gnd OAI21X1_280/C vdd NAND2X1
XNAND2X1_369 BUFX4_75/Y OAI21X1_401/B gnd OAI21X1_372/C vdd NAND2X1
XNAND2X1_358 BUFX4_122/Y OAI21X1_349/Y gnd OAI21X1_350/C vdd NAND2X1
XNAND2X1_347 BUFX4_20/Y MUX2X1_2/Y gnd NOR2X1_170/B vdd NAND2X1
XNOR2X1_391 BUFX2_63/A BUFX2_64/A gnd NOR2X1_391/Y vdd NOR2X1
XNOR2X1_380 NOR2X1_380/A NOR2X1_380/B gnd NOR2X1_380/Y vdd NOR2X1
XFILL_25_3_0 gnd vdd FILL
XFILL_0_3_0 gnd vdd FILL
XINVX4_6 operand_A[17] gnd INVX4_6/Y vdd INVX4
XOAI21X1_875 OAI21X1_875/A NOR2X1_87/B NOR2X1_22/A gnd OAI22X1_29/B vdd OAI21X1
XOAI21X1_886 OAI21X1_2/C OAI21X1_901/A OAI21X1_886/C gnd OAI21X1_886/Y vdd OAI21X1
XOAI21X1_897 BUFX4_65/Y OAI21X1_4/C BUFX4_100/Y gnd NOR2X1_495/A vdd OAI21X1
XOAI21X1_831 NOR2X1_463/Y OAI21X1_17/Y NAND2X1_40/B gnd INVX1_309/A vdd OAI21X1
XOAI21X1_820 BUFX4_65/Y INVX1_307/Y OAI21X1_820/C gnd NOR2X1_460/B vdd OAI21X1
XOAI21X1_842 OAI21X1_842/A OAI21X1_842/B BUFX4_100/Y gnd OAI21X1_843/C vdd OAI21X1
XOAI21X1_864 NOR2X1_485/B OAI21X1_7/C BUFX4_138/Y gnd OAI21X1_864/Y vdd OAI21X1
XOAI21X1_853 NOR2X1_473/Y OAI21X1_853/B INVX8_10/A gnd AND2X2_65/A vdd OAI21X1
XFILL_8_4_0 gnd vdd FILL
XFILL_16_3_0 gnd vdd FILL
XNAND3X1_9 NAND3X1_9/A NAND3X1_9/B OR2X2_9/Y gnd NAND3X1_9/Y vdd NAND3X1
XOAI21X1_149 NOR2X1_97/A INVX1_76/Y AND2X2_6/Y gnd OAI21X1_150/A vdd OAI21X1
XOAI21X1_105 INVX2_2/Y MUX2X1_1/S OAI21X1_105/C gnd INVX1_63/A vdd OAI21X1
XOAI21X1_138 BUFX4_190/Y MUX2X1_18/Y OAI21X1_138/C gnd OAI21X1_265/B vdd OAI21X1
XOAI21X1_127 BUFX4_192/Y MUX2X1_14/Y OAI21X1_127/C gnd MUX2X1_30/B vdd OAI21X1
XBUFX2_3 BUFX2_3/A gnd result[0] vdd BUFX2
XOAI21X1_116 INVX2_24/Y MUX2X1_5/S OAI21X1_116/C gnd OAI21X1_211/B vdd OAI21X1
XNAND2X1_133 BUFX4_46/Y operand_A[41] gnd OAI21X1_82/C vdd NAND2X1
XNAND2X1_122 MUX2X1_5/S operand_A[47] gnd OAI21X1_71/C vdd NAND2X1
XNAND2X1_111 NOR2X1_82/A MUX2X1_5/Y gnd OAI21X1_62/C vdd NAND2X1
XNAND2X1_177 MUX2X1_51/S MUX2X1_30/A gnd OAI21X1_133/C vdd NAND2X1
XNAND2X1_100 BUFX4_66/Y MUX2X1_1/Y gnd OAI21X1_51/C vdd NAND2X1
XNAND2X1_155 BUFX4_53/Y operand_A[2] gnd OAI21X1_111/C vdd NAND2X1
XNAND2X1_166 BUFX4_20/Y INVX1_149/A gnd OAI21X1_122/C vdd NAND2X1
XNAND2X1_144 MUX2X1_8/S operand_A[22] gnd OAI21X1_99/C vdd NAND2X1
XNAND2X1_188 BUFX4_21/Y MUX2X1_20/Y gnd OAI21X1_145/C vdd NAND2X1
XNAND2X1_199 operand_A[2] NOR2X1_19/B gnd OAI21X1_743/C vdd NAND2X1
XOAI21X1_650 operand_B[21] INVX4_4/Y OAI21X1_650/C gnd OAI21X1_650/Y vdd OAI21X1
XINVX2_3 operand_B[20] gnd INVX2_3/Y vdd INVX2
XOAI21X1_661 INVX1_219/A OAI21X1_661/B OAI21X1_661/C gnd OAI21X1_661/Y vdd OAI21X1
XOAI21X1_672 INVX1_162/A OAI21X1_672/B OAI21X1_672/C gnd OAI21X1_672/Y vdd OAI21X1
XOAI21X1_683 INVX2_22/Y MUX2X1_3/S OAI21X1_55/C gnd OAI21X1_683/Y vdd OAI21X1
XOAI21X1_694 MUX2X1_64/S MUX2X1_75/Y NAND3X1_56/Y gnd OAI21X1_695/B vdd OAI21X1
XAOI21X1_3 NOR2X1_10/Y XOR2X1_2/Y NOR2X1_9/Y gnd OAI21X1_3/C vdd AOI21X1
XXNOR2X1_33 XNOR2X1_33/A INVX1_148/A gnd XNOR2X1_33/Y vdd XNOR2X1
XXNOR2X1_11 operand_A[23] operand_B[23] gnd XNOR2X1_46/B vdd XNOR2X1
XINVX1_90 INVX1_90/A gnd INVX1_90/Y vdd INVX1
XXNOR2X1_44 XNOR2X1_44/A OAI21X1_2/C gnd XNOR2X1_44/Y vdd XNOR2X1
XXNOR2X1_22 operand_A[15] operand_B[15] gnd XNOR2X1_22/Y vdd XNOR2X1
XBUFX2_10 BUFX2_10/A gnd result[7] vdd BUFX2
XBUFX2_43 BUFX2_43/A gnd result[40] vdd BUFX2
XBUFX2_65 BUFX2_65/A gnd result[62] vdd BUFX2
XBUFX2_54 BUFX2_54/A gnd result[51] vdd BUFX2
XBUFX2_32 BUFX2_32/A gnd result[29] vdd BUFX2
XFILL_31_1_0 gnd vdd FILL
XBUFX2_21 BUFX2_21/A gnd result[18] vdd BUFX2
XNOR2X1_1 INVX2_1/Y INVX2_2/Y gnd NOR2X1_1/Y vdd NOR2X1
XFILL_22_1_0 gnd vdd FILL
XAOI21X1_44 AOI21X1_44/A OAI21X1_93/Y NOR2X1_93/Y gnd AOI21X1_44/Y vdd AOI21X1
XAOI21X1_99 OR2X2_12/B OR2X2_12/A BUFX4_93/Y gnd AOI22X1_9/D vdd AOI21X1
XAOI21X1_77 INVX2_62/A NOR2X1_144/Y BUFX4_29/Y gnd AOI21X1_77/Y vdd AOI21X1
XAOI21X1_33 NAND2X1_55/B NOR2X1_69/Y NOR2X1_68/Y gnd INVX1_32/A vdd AOI21X1
XAOI21X1_88 INVX8_18/A INVX1_296/A OAI22X1_5/Y gnd NAND3X1_12/B vdd AOI21X1
XOAI21X1_6 NOR2X1_6/B OAI21X1_6/B OAI21X1_6/C gnd OAI21X1_6/Y vdd OAI21X1
XAOI21X1_66 OR2X2_7/Y AOI21X1_66/B BUFX4_172/Y gnd AOI21X1_66/Y vdd AOI21X1
XAOI21X1_55 AND2X2_10/Y AOI21X1_55/B AOI21X1_55/C gnd NOR2X1_485/B vdd AOI21X1
XAOI21X1_22 INVX1_279/A NAND2X1_68/Y NOR2X1_54/Y gnd OAI21X1_28/B vdd AOI21X1
XAOI21X1_11 NAND2X1_42/Y NOR2X1_35/Y NOR2X1_34/Y gnd OAI21X1_17/C vdd AOI21X1
XFILL_5_2_0 gnd vdd FILL
XFILL_13_1_0 gnd vdd FILL
XOAI22X1_30 BUFX4_78/Y OAI22X1_30/B OAI22X1_30/C OAI22X1_30/D gnd OAI22X1_30/Y vdd
+ OAI22X1
XOAI21X1_491 INVX2_52/Y MUX2X1_7/S OAI21X1_491/C gnd INVX1_205/A vdd OAI21X1
XOAI21X1_480 INVX1_188/Y BUFX4_73/Y OAI21X1_480/C gnd INVX1_217/A vdd OAI21X1
XBUFX4_149 NOR2X1_89/Y gnd BUFX4_149/Y vdd BUFX4
XNOR2X1_209 INVX2_73/Y INVX1_173/Y gnd NOR2X1_210/B vdd NOR2X1
XBUFX4_138 NOR2X1_72/Y gnd BUFX4_138/Y vdd BUFX4
XBUFX4_127 INVX8_3/Y gnd MUX2X1_27/S vdd BUFX4
XBUFX4_116 operand_B[5] gnd BUFX4_116/Y vdd BUFX4
XBUFX4_105 NOR2X1_45/Y gnd BUFX4_105/Y vdd BUFX4
XINVX1_330 reset gnd DFFSR_1/R vdd INVX1
XFILL_20_4_1 gnd vdd FILL
XAOI21X1_389 INVX2_94/Y BUFX4_60/Y NAND2X1_640/Y gnd NAND2X1_641/B vdd AOI21X1
XAOI21X1_345 NOR2X1_37/Y BUFX4_150/Y AOI21X1_345/C gnd OAI21X1_835/C vdd AOI21X1
XAOI21X1_312 XNOR2X1_17/Y OAI21X1_744/B BUFX4_92/Y gnd OAI21X1_744/C vdd AOI21X1
XAOI21X1_301 XOR2X1_3/Y INVX8_14/A OAI21X1_702/Y gnd NAND2X1_567/B vdd AOI21X1
XAOI21X1_323 XNOR2X1_19/Y OAI21X1_781/A OAI21X1_779/Y gnd AOI21X1_324/C vdd AOI21X1
XAOI21X1_356 BUFX4_85/Y NOR2X1_474/Y OAI21X1_855/Y gnd AND2X2_65/B vdd AOI21X1
XAOI21X1_334 XNOR2X1_7/Y INVX2_93/Y BUFX4_31/Y gnd OAI21X1_812/C vdd AOI21X1
XDFFPOSX1_11 BUFX2_13/A CLKBUF1_2/Y AOI22X1_40/Y gnd vdd DFFPOSX1
XAOI21X1_367 BUFX4_77/Y MUX2X1_123/Y INVX8_9/Y gnd OAI22X1_28/C vdd AOI21X1
XAOI21X1_378 BUFX4_138/Y XNOR2X1_43/Y NAND2X1_631/Y gnd AOI22X1_49/C vdd AOI21X1
XDFFPOSX1_55 OR2X2_37/A CLKBUF1_5/Y DFFPOSX1_55/D gnd vdd DFFPOSX1
XDFFPOSX1_44 BUFX2_46/A CLKBUF1_8/Y DFFPOSX1_44/D gnd vdd DFFPOSX1
XDFFPOSX1_33 BUFX2_35/A CLKBUF1_8/Y AOI21X1_65/Y gnd vdd DFFPOSX1
XDFFPOSX1_22 OR2X2_48/B DFFSR_1/CLK AND2X2_72/Y gnd vdd DFFPOSX1
XFILL_28_5_1 gnd vdd FILL
XFILL_27_0_0 gnd vdd FILL
XFILL_2_0_0 gnd vdd FILL
XFILL_3_5_1 gnd vdd FILL
XFILL_11_4_1 gnd vdd FILL
XFILL_19_5_1 gnd vdd FILL
XFILL_18_0_0 gnd vdd FILL
XNAND2X1_507 INVX2_84/A OAI21X1_583/B gnd OAI21X1_590/C vdd NAND2X1
XINVX1_171 INVX1_171/A gnd INVX1_171/Y vdd INVX1
XINVX1_182 INVX1_182/A gnd INVX1_182/Y vdd INVX1
XNAND2X1_518 BUFX4_70/Y INVX1_254/Y gnd OAI21X1_614/C vdd NAND2X1
XINVX1_160 INVX1_160/A gnd INVX1_160/Y vdd INVX1
XINVX1_193 INVX1_193/A gnd INVX1_193/Y vdd INVX1
XNAND2X1_529 NOR2X1_376/Y NOR2X1_377/Y gnd NOR2X1_380/A vdd NAND2X1
XAOI21X1_186 INVX1_212/Y NOR2X1_273/Y BUFX4_30/Y gnd OAI21X1_509/C vdd AOI21X1
XAOI21X1_175 INVX1_201/A INVX1_204/A NOR2X1_258/B gnd INVX1_208/A vdd AOI21X1
XAOI21X1_197 BUFX4_143/Y XNOR2X1_39/Y NAND3X1_32/Y gnd AOI21X1_198/B vdd AOI21X1
XAOI21X1_131 OAI21X1_393/Y AOI21X1_131/B NOR2X1_207/Y gnd DFFPOSX1_43/D vdd AOI21X1
XAOI21X1_164 NAND2X1_427/B NOR2X1_231/B INVX1_194/Y gnd NAND3X1_29/B vdd AOI21X1
XAOI21X1_153 NOR2X1_232/Y INVX4_21/A NOR2X1_233/Y gnd NOR2X1_249/B vdd AOI21X1
XAOI21X1_142 INVX1_250/A INVX1_176/Y BUFX4_159/Y gnd OR2X2_44/B vdd AOI21X1
XAOI21X1_120 INVX4_18/A NOR2X1_195/Y OR2X2_18/Y gnd NAND3X1_18/B vdd AOI21X1
XFILL_20_2 gnd vdd FILL
XBUFX4_7 BUFX4_9/A gnd BUFX4_7/Y vdd BUFX4
XOAI21X1_309 INVX1_134/Y MUX2X1_71/S OAI21X1_309/C gnd OAI21X1_847/A vdd OAI21X1
XNAND2X1_348 BUFX4_75/Y INVX1_159/A gnd OAI21X1_337/C vdd NAND2X1
XNAND2X1_315 BUFX4_114/Y OAI22X1_27/A gnd NAND3X1_12/A vdd NAND2X1
XNAND2X1_337 BUFX4_120/Y OAI21X1_323/Y gnd OAI21X1_324/C vdd NAND2X1
XNAND2X1_326 MUX2X1_71/S MUX2X1_27/B gnd OAI21X1_309/C vdd NAND2X1
XNAND2X1_304 BUFX4_20/Y OAI21X1_411/B gnd OAI21X1_281/C vdd NAND2X1
XNAND2X1_359 BUFX4_23/Y INVX1_196/A gnd OAI21X1_351/C vdd NAND2X1
XFILL_25_3_1 gnd vdd FILL
XNOR2X1_381 BUFX2_42/A BUFX2_43/A gnd NOR2X1_381/Y vdd NOR2X1
XNOR2X1_392 BUFX2_61/A BUFX2_62/A gnd NOR2X1_392/Y vdd NOR2X1
XNOR2X1_370 operand_A[63] operand_B[63] gnd NOR2X1_371/A vdd NOR2X1
XINVX4_7 operand_A[4] gnd INVX4_7/Y vdd INVX4
XFILL_0_3_1 gnd vdd FILL
XOAI21X1_832 INVX2_93/Y OAI21X1_17/A OAI21X1_17/C gnd OAI21X1_833/A vdd OAI21X1
XOAI21X1_821 BUFX4_155/Y XNOR2X1_7/Y OR2X2_48/A gnd NOR2X1_460/A vdd OAI21X1
XOAI21X1_810 NOR2X1_198/B BUFX4_77/Y OAI21X1_810/C gnd AOI22X1_38/D vdd OAI21X1
XOAI21X1_898 AND2X2_71/Y OAI21X1_898/B OAI21X1_898/C gnd AND2X2_72/A vdd OAI21X1
XOAI21X1_887 INVX1_320/Y NOR2X1_80/A OAI21X1_887/C gnd AOI22X1_50/C vdd OAI21X1
XOAI21X1_854 operand_B[14] operand_A[14] BUFX4_1/Y gnd OAI21X1_855/C vdd OAI21X1
XOAI21X1_843 BUFX4_100/Y INVX1_308/Y OAI21X1_843/C gnd OAI21X1_843/Y vdd OAI21X1
XOAI21X1_865 operand_B[16] operand_A[16] BUFX4_1/Y gnd AND2X2_66/A vdd OAI21X1
XOAI21X1_876 operand_A[18] operand_B[18] BUFX4_3/Y gnd OAI21X1_877/C vdd OAI21X1
XFILL_8_4_1 gnd vdd FILL
XFILL_16_3_1 gnd vdd FILL
XOAI21X1_106 INVX2_50/Y MUX2X1_6/S OAI21X1_106/C gnd OAI21X1_106/Y vdd OAI21X1
XOAI21X1_128 BUFX4_131/Y MUX2X1_30/B OAI21X1_128/C gnd NOR2X1_177/B vdd OAI21X1
XOAI21X1_117 BUFX4_190/Y MUX2X1_12/Y OAI21X1_117/C gnd INVX1_67/A vdd OAI21X1
XOAI21X1_139 INVX1_70/Y MUX2X1_87/S OAI21X1_139/C gnd MUX2X1_36/A vdd OAI21X1
XBUFX2_4 BUFX2_4/A gnd result[1] vdd BUFX2
XNAND2X1_178 MUX2X1_7/S operand_A[42] gnd OAI21X1_412/C vdd NAND2X1
XNAND2X1_112 BUFX4_48/Y operand_A[59] gnd OAI21X1_61/C vdd NAND2X1
XNAND2X1_123 BUFX4_68/Y INVX1_87/A gnd OAI21X1_72/C vdd NAND2X1
XNAND2X1_167 MUX2X1_7/S operand_A[62] gnd OAI21X1_628/A vdd NAND2X1
XNAND2X1_134 MUX2X1_97/S OAI21X1_82/Y gnd OAI21X1_83/C vdd NAND2X1
XNAND2X1_189 INVX2_49/A AND2X2_7/Y gnd INVX1_74/A vdd NAND2X1
XNAND2X1_101 BUFX4_50/Y operand_A[3] gnd OAI21X1_52/C vdd NAND2X1
XNAND2X1_156 BUFX4_66/Y INVX1_65/Y gnd OAI21X1_112/C vdd NAND2X1
XNAND2X1_145 BUFX4_76/Y OAI21X1_99/Y gnd OAI21X1_100/C vdd NAND2X1
XOAI21X1_662 AOI22X1_30/Y NOR2X1_312/A OAI21X1_662/C gnd AND2X2_49/A vdd OAI21X1
XOAI21X1_673 NOR2X1_423/Y OR2X2_29/B OAI21X1_673/C gnd OAI21X1_673/Y vdd OAI21X1
XOAI21X1_651 OAI21X1_651/A OAI21X1_651/B NOR2X1_120/Y gnd NAND3X1_54/C vdd OAI21X1
XAOI21X1_4 AOI21X1_4/A OR2X2_49/B NOR2X1_11/Y gnd OAI21X1_6/C vdd AOI21X1
XOAI21X1_684 INVX1_286/Y INVX8_1/A OAI21X1_684/C gnd INVX1_287/A vdd OAI21X1
XOAI21X1_640 OAI21X1_640/A NOR2X1_60/A OAI21X1_640/C gnd AOI22X1_29/C vdd OAI21X1
XINVX2_4 operand_A[20] gnd INVX2_4/Y vdd INVX2
XXNOR2X1_12 operand_B[21] operand_A[21] gnd AND2X2_71/B vdd XNOR2X1
XXNOR2X1_23 operand_B[14] operand_A[14] gnd XNOR2X1_23/Y vdd XNOR2X1
XOAI21X1_695 NOR2X1_22/A OAI21X1_695/B OAI21X1_695/C gnd OAI21X1_695/Y vdd OAI21X1
XBUFX2_33 BUFX2_33/A gnd result[30] vdd BUFX2
XBUFX2_44 OR2X2_36/B gnd result[41] vdd BUFX2
XXNOR2X1_34 XNOR2X1_34/A INVX4_21/Y gnd XNOR2X1_34/Y vdd XNOR2X1
XXNOR2X1_45 XNOR2X1_45/A AND2X2_71/B gnd XNOR2X1_45/Y vdd XNOR2X1
XINVX1_80 INVX1_80/A gnd INVX1_80/Y vdd INVX1
XINVX1_91 INVX1_91/A gnd INVX1_91/Y vdd INVX1
XBUFX2_11 BUFX2_11/A gnd result[8] vdd BUFX2
XBUFX2_22 BUFX2_22/A gnd result[19] vdd BUFX2
XBUFX2_66 BUFX2_66/A gnd result[63] vdd BUFX2
XBUFX2_55 BUFX2_55/A gnd result[52] vdd BUFX2
XFILL_31_1_1 gnd vdd FILL
XNOR2X1_2 INVX1_1/Y INVX4_2/Y gnd NOR2X1_2/Y vdd NOR2X1
XAOI21X1_34 INVX1_34/Y OAI21X1_34/Y AND2X2_2/Y gnd NOR2X1_96/B vdd AOI21X1
XFILL_22_1_1 gnd vdd FILL
XAOI21X1_23 INVX1_280/A OAI21X1_8/A INVX1_80/A gnd OAI21X1_28/C vdd AOI21X1
XAOI21X1_12 NOR2X1_37/Y INVX1_21/Y NOR2X1_36/Y gnd INVX1_312/A vdd AOI21X1
XAOI21X1_89 INVX4_19/A INVX2_64/A INVX2_63/Y gnd AOI21X1_90/B vdd AOI21X1
XAOI21X1_56 AND2X2_2/Y NOR2X1_119/Y AOI21X1_56/C gnd AOI21X1_56/Y vdd AOI21X1
XAOI21X1_45 AND2X2_5/Y AND2X2_6/A INVX1_75/Y gnd AOI21X1_45/Y vdd AOI21X1
XAOI21X1_67 INVX4_20/A AND2X2_52/A OR2X2_8/Y gnd NAND3X1_8/B vdd AOI21X1
XAOI21X1_78 BUFX4_186/Y AOI21X1_78/B NOR2X1_145/Y gnd NOR2X1_435/B vdd AOI21X1
XOAI21X1_7 INVX1_11/Y OAI21X1_7/B OAI21X1_7/C gnd OAI21X1_7/Y vdd OAI21X1
XFILL_5_2_1 gnd vdd FILL
XOAI22X1_20 BUFX4_64/Y INVX1_251/Y BUFX4_157/Y INVX2_88/Y gnd OAI22X1_20/Y vdd OAI22X1
XFILL_13_1_1 gnd vdd FILL
XOAI22X1_31 OAI22X1_31/A OAI22X1_31/B OAI22X1_31/C OAI22X1_31/D gnd OAI22X1_31/Y vdd
+ OAI22X1
XOAI21X1_492 INVX1_205/Y MUX2X1_98/S OAI21X1_492/C gnd INVX1_206/A vdd OAI21X1
XOAI21X1_481 INVX1_178/Y MUX2X1_66/S OAI21X1_481/C gnd MUX2X1_54/A vdd OAI21X1
XOAI21X1_470 INVX1_196/Y BUFX4_25/Y OAI21X1_470/C gnd OAI22X1_23/C vdd OAI21X1
XBUFX4_139 NOR2X1_72/Y gnd INVX8_11/A vdd BUFX4
XBUFX4_106 NOR2X1_45/Y gnd INVX8_6/A vdd BUFX4
XBUFX4_117 INVX8_3/Y gnd MUX2X1_2/S vdd BUFX4
XBUFX4_128 operand_B[2] gnd INVX8_3/A vdd BUFX4
XINVX1_320 MUX2X1_33/Y gnd INVX1_320/Y vdd INVX1
XFILL_1_1 gnd vdd FILL
XDFFPOSX1_34 BUFX2_36/A CLKBUF1_3/Y AOI21X1_69/Y gnd vdd DFFPOSX1
XDFFPOSX1_45 BUFX2_47/A CLKBUF1_8/Y DFFPOSX1_45/D gnd vdd DFFPOSX1
XDFFPOSX1_23 BUFX2_25/A CLKBUF1_1/Y OAI21X1_905/Y gnd vdd DFFPOSX1
XAOI21X1_335 INVX8_10/A INVX1_172/Y BUFX4_80/Y gnd OAI21X1_813/C vdd AOI21X1
XAOI21X1_379 AND2X2_1/B INVX1_315/A OAI21X1_3/Y gnd XNOR2X1_44/A vdd AOI21X1
XAOI21X1_313 NOR2X1_16/Y BUFX4_150/Y BUFX4_14/Y gnd NAND2X1_594/A vdd AOI21X1
XDFFPOSX1_12 BUFX2_14/A CLKBUF1_2/Y AOI22X1_42/Y gnd vdd DFFPOSX1
XAOI21X1_324 INVX8_10/A OAI21X1_780/Y AOI21X1_324/C gnd AOI21X1_325/B vdd AOI21X1
XAOI21X1_302 BUFX4_86/Y NOR2X1_427/Y NAND2X1_567/Y gnd AND2X2_53/B vdd AOI21X1
XAOI21X1_368 INVX4_26/Y OR2X2_46/Y BUFX4_31/Y gnd OAI21X1_868/C vdd AOI21X1
XAOI21X1_357 BUFX4_114/Y INVX1_189/Y OAI21X1_853/B gnd NOR2X1_475/B vdd AOI21X1
XAOI21X1_346 INVX8_4/A OR2X2_44/Y NOR2X1_466/Y gnd OAI21X1_841/B vdd AOI21X1
XDFFPOSX1_56 BUFX2_58/A CLKBUF1_4/Y DFFPOSX1_56/D gnd vdd DFFPOSX1
XFILL_27_0_1 gnd vdd FILL
XFILL_2_0_1 gnd vdd FILL
XFILL_18_0_1 gnd vdd FILL
XINVX1_161 operand_B[41] gnd INVX1_161/Y vdd INVX1
XINVX1_194 INVX1_194/A gnd INVX1_194/Y vdd INVX1
XINVX1_172 INVX1_172/A gnd INVX1_172/Y vdd INVX1
XNAND2X1_519 INVX4_18/A MUX2X1_64/Y gnd NAND3X1_36/A vdd NAND2X1
XNAND2X1_508 BUFX4_186/Y NOR2X1_212/B gnd NAND2X1_508/Y vdd NAND2X1
XINVX1_183 INVX1_183/A gnd INVX1_183/Y vdd INVX1
XINVX1_150 INVX1_150/A gnd INVX1_150/Y vdd INVX1
XAOI21X1_110 AOI21X1_110/A OAI21X1_347/Y NOR2X1_172/Y gnd DFFPOSX1_40/D vdd AOI21X1
XAOI21X1_132 INVX2_74/A OAI21X1_409/B BUFX4_28/Y gnd OAI21X1_409/C vdd AOI21X1
XAOI21X1_121 OR2X2_7/B OAI21X1_391/Y AND2X2_18/Y gnd NOR2X1_196/B vdd AOI21X1
XAOI21X1_198 OAI21X1_531/Y AOI21X1_198/B NOR2X1_289/Y gnd DFFPOSX1_54/D vdd AOI21X1
XAOI21X1_176 INVX1_207/Y AND2X2_26/A INVX1_208/Y gnd NOR2X1_272/B vdd AOI21X1
XAOI21X1_165 INVX1_153/A INVX1_198/Y NAND3X1_29/Y gnd OAI21X1_472/C vdd AOI21X1
XAOI21X1_143 OR2X2_7/B INVX1_176/A OR2X2_44/A gnd NOR2X1_467/B vdd AOI21X1
XAOI21X1_154 BUFX4_179/Y INVX1_56/A NOR2X1_235/Y gnd OR2X2_25/A vdd AOI21X1
XAOI21X1_187 BUFX4_164/Y INVX1_119/Y INVX4_11/A gnd OAI21X1_515/A vdd AOI21X1
XBUFX4_8 BUFX4_9/A gnd BUFX4_8/Y vdd BUFX4
XNAND2X1_316 MUX2X1_99/S OAI21X1_176/Y gnd OAI21X1_299/C vdd NAND2X1
XNAND2X1_349 BUFX4_120/Y OAI21X1_337/Y gnd OAI21X1_338/C vdd NAND2X1
XNAND2X1_305 AOI22X1_7/Y NOR2X1_149/Y gnd AOI21X1_80/C vdd NAND2X1
XNAND2X1_338 BUFX4_23/Y OAI21X1_443/B gnd OAI21X1_325/C vdd NAND2X1
XNAND2X1_327 BUFX4_22/Y OAI21X1_847/A gnd OAI21X1_310/C vdd NAND2X1
XNOR2X1_360 OR2X2_43/B MUX2X1_63/Y gnd NOR2X1_360/Y vdd NOR2X1
XNOR2X1_393 OR2X2_37/Y NOR2X1_393/B gnd NOR2X1_393/Y vdd NOR2X1
XNOR2X1_382 BUFX2_47/A BUFX2_48/A gnd NOR2X1_382/Y vdd NOR2X1
XNOR2X1_371 NOR2X1_371/A AND2X2_44/Y gnd INVX4_25/A vdd NOR2X1
XINVX4_8 operand_A[25] gnd INVX4_8/Y vdd INVX4
XOAI21X1_844 INVX1_309/Y NOR2X1_37/Y XNOR2X1_41/B gnd NAND3X1_65/C vdd OAI21X1
XOAI21X1_833 OAI21X1_833/A NAND2X1_40/B BUFX4_105/Y gnd OAI21X1_835/A vdd OAI21X1
XOAI21X1_811 INVX1_306/Y INVX2_17/A OAI21X1_17/B gnd INVX2_93/A vdd OAI21X1
XOAI21X1_822 OAI21X1_822/A NOR2X1_459/Y NOR2X1_460/Y gnd OAI21X1_822/Y vdd OAI21X1
XOAI21X1_855 BUFX4_65/Y OAI21X1_855/B OAI21X1_855/C gnd OAI21X1_855/Y vdd OAI21X1
XOAI21X1_800 AND2X2_57/Y OAI21X1_800/B INVX8_10/A gnd OAI21X1_801/C vdd OAI21X1
XOAI21X1_866 XNOR2X1_25/Y BUFX4_155/Y AND2X2_66/Y gnd NOR2X1_483/A vdd OAI21X1
XOAI21X1_888 OAI22X1_12/B BUFX4_171/Y BUFX4_111/Y gnd OAI21X1_888/Y vdd OAI21X1
XOAI21X1_899 XNOR2X1_44/A NOR2X1_6/A OAI21X1_6/B gnd AND2X2_73/A vdd OAI21X1
XOAI21X1_877 BUFX4_65/Y INVX1_317/Y OAI21X1_877/C gnd NOR2X1_488/B vdd OAI21X1
XOAI21X1_129 INVX2_52/Y MUX2X1_5/S OAI21X1_511/C gnd OAI21X1_129/Y vdd OAI21X1
XOAI21X1_107 INVX1_63/Y BUFX4_68/Y OAI21X1_107/C gnd OAI21X1_107/Y vdd OAI21X1
XOAI21X1_118 INVX2_20/Y MUX2X1_1/S OAI21X1_118/C gnd INVX1_68/A vdd OAI21X1
XBUFX2_5 BUFX2_5/A gnd result[2] vdd BUFX2
XNAND2X1_179 INVX8_1/A OAI21X1_135/Y gnd OAI21X1_136/C vdd NAND2X1
XNAND2X1_168 BUFX4_70/Y MUX2X1_13/Y gnd OAI21X1_125/C vdd NAND2X1
XNAND2X1_135 MUX2X1_71/S OAI21X1_83/Y gnd OAI21X1_84/C vdd NAND2X1
XNAND2X1_124 MUX2X1_30/S OAI21X1_72/Y gnd OAI21X1_73/C vdd NAND2X1
XNAND2X1_113 BUFX4_133/Y OAI21X1_62/Y gnd OAI21X1_66/C vdd NAND2X1
XNAND2X1_157 BUFX4_43/Y operand_A[4] gnd OAI21X1_113/C vdd NAND2X1
XNAND2X1_102 MUX2X1_7/S operand_A[5] gnd OAI21X1_53/C vdd NAND2X1
XNAND2X1_146 BUFX4_119/Y OAI21X1_100/Y gnd OAI21X1_101/C vdd NAND2X1
XNOR2X1_190 NOR2X1_190/A NOR2X1_190/B gnd INVX1_162/A vdd NOR2X1
XOAI21X1_663 AND2X2_49/Y OAI21X1_663/B INVX2_89/Y gnd OAI21X1_663/Y vdd OAI21X1
XOAI21X1_674 OAI21X1_674/A NOR2X1_412/B AND2X2_50/Y gnd NOR2X1_424/B vdd OAI21X1
XOAI21X1_652 NAND2X1_59/A NAND2X1_58/B NAND2X1_55/B gnd NAND3X1_53/B vdd OAI21X1
XOAI21X1_630 OAI21X1_630/A MUX2X1_62/S OAI21X1_630/C gnd NOR2X1_373/B vdd OAI21X1
XAOI21X1_5 NOR2X1_6/Y OAI21X1_3/Y OAI21X1_6/Y gnd INVX1_10/A vdd AOI21X1
XOAI21X1_685 INVX2_21/Y BUFX4_43/Y OAI21X1_685/C gnd INVX1_288/A vdd OAI21X1
XOAI21X1_641 XNOR2X1_41/B NAND2X1_39/B NAND2X1_36/B gnd AOI22X1_29/B vdd OAI21X1
XOAI21X1_696 INVX8_14/A NOR2X1_426/Y NOR2X1_410/B gnd AND2X2_51/B vdd OAI21X1
XINVX2_5 operand_B[18] gnd INVX2_5/Y vdd INVX2
XXNOR2X1_35 XNOR2X1_35/A INVX4_22/Y gnd XNOR2X1_35/Y vdd XNOR2X1
XXNOR2X1_46 OR2X2_49/Y XNOR2X1_46/B gnd XNOR2X1_46/Y vdd XNOR2X1
XXNOR2X1_13 operand_B[20] operand_A[20] gnd XNOR2X1_13/Y vdd XNOR2X1
XXNOR2X1_24 operand_B[17] operand_A[17] gnd INVX4_26/A vdd XNOR2X1
XBUFX2_34 BUFX2_34/A gnd result[31] vdd BUFX2
XBUFX2_45 BUFX2_45/A gnd result[42] vdd BUFX2
XBUFX2_56 BUFX2_56/A gnd result[53] vdd BUFX2
XBUFX2_23 BUFX2_23/A gnd result[20] vdd BUFX2
XBUFX2_67 BUFX2_67/A gnd zero_flag vdd BUFX2
XINVX1_70 INVX1_70/A gnd INVX1_70/Y vdd INVX1
XINVX1_81 INVX1_81/A gnd INVX1_81/Y vdd INVX1
XBUFX2_12 BUFX2_12/A gnd result[9] vdd BUFX2
XINVX1_92 INVX1_92/A gnd INVX1_92/Y vdd INVX1
XNOR2X1_3 NOR2X1_3/A NOR2X1_3/B gnd NOR2X1_3/Y vdd NOR2X1
XAOI21X1_35 INVX4_1/Y NOR2X1_96/B OAI21X1_35/Y gnd NOR2X1_91/A vdd AOI21X1
XAOI21X1_46 AND2X2_9/Y INVX1_25/A AOI21X1_46/C gnd AOI21X1_46/Y vdd AOI21X1
XAOI21X1_68 NAND3X1_9/A XNOR2X1_30/Y NAND3X1_8/Y gnd AOI21X1_69/B vdd AOI21X1
XAOI21X1_57 NOR2X1_120/Y NAND2X1_66/Y AOI21X1_57/C gnd AOI21X1_57/Y vdd AOI21X1
XAOI21X1_24 NAND2X1_73/Y NOR2X1_57/Y NOR2X1_22/Y gnd OAI21X1_29/B vdd AOI21X1
XAOI21X1_13 NAND2X1_43/Y NOR2X1_40/Y NOR2X1_39/Y gnd OAI21X1_18/C vdd AOI21X1
XAOI21X1_79 BUFX4_41/Y AND2X2_20/A NOR2X1_150/Y gnd INVX1_119/A vdd AOI21X1
XOAI21X1_8 OAI21X1_8/A OAI21X1_8/B XOR2X1_4/Y gnd OAI21X1_9/B vdd OAI21X1
XOAI22X1_32 OAI22X1_32/A OAI22X1_32/B OAI22X1_32/C OAI22X1_32/D gnd OAI22X1_32/Y vdd
+ OAI22X1
XOAI22X1_21 OAI22X1_21/A OAI22X1_21/B OAI22X1_2/D BUFX4_81/Y gnd OAI22X1_21/Y vdd
+ OAI22X1
XOAI22X1_10 OAI22X1_1/B OR2X2_10/A INVX1_124/Y INVX8_8/Y gnd OAI22X1_30/D vdd OAI22X1
XOAI21X1_493 INVX1_206/Y BUFX4_131/Y OAI21X1_493/C gnd MUX2X1_55/A vdd OAI21X1
XOAI21X1_471 OAI22X1_23/C MUX2X1_57/S BUFX4_84/Y gnd OAI22X1_8/D vdd OAI21X1
XOAI21X1_482 INVX1_160/Y BUFX4_18/Y OAI21X1_482/C gnd MUX2X1_42/A vdd OAI21X1
XOAI21X1_460 OAI21X1_460/A NOR2X1_22/A OAI21X1_460/C gnd NAND3X1_25/A vdd OAI21X1
XFILL_32_4_0 gnd vdd FILL
XFILL_23_4_0 gnd vdd FILL
XBUFX4_107 NOR2X1_45/Y gnd BUFX4_107/Y vdd BUFX4
XBUFX4_118 INVX8_3/Y gnd MUX2X1_30/S vdd BUFX4
XFILL_6_5_0 gnd vdd FILL
XFILL_14_4_0 gnd vdd FILL
XBUFX4_129 operand_B[2] gnd NOR2X1_83/A vdd BUFX4
XINVX1_321 INVX1_321/A gnd INVX1_321/Y vdd INVX1
XOAI21X1_290 MUX2X1_2/S OAI21X1_290/B OAI21X1_290/C gnd MUX2X1_31/B vdd OAI21X1
XINVX1_310 INVX1_310/A gnd INVX1_310/Y vdd INVX1
XFILL_1_2 gnd vdd FILL
XAOI21X1_303 NAND2X1_571/Y NAND2X1_575/Y BUFX4_162/Y gnd OAI21X1_714/A vdd AOI21X1
XAOI21X1_314 NOR2X1_438/Y OAI21X1_732/Y NOR2X1_434/Y gnd DFFPOSX1_4/D vdd AOI21X1
XAOI21X1_325 AOI21X1_325/A AOI21X1_325/B NOR2X1_445/Y gnd DFFPOSX1_7/D vdd AOI21X1
XDFFPOSX1_35 BUFX2_37/A CLKBUF1_3/Y AOI21X1_76/Y gnd vdd DFFPOSX1
XDFFPOSX1_57 BUFX2_59/A CLKBUF1_4/Y DFFPOSX1_57/D gnd vdd DFFPOSX1
XDFFPOSX1_46 BUFX2_48/A DFFSR_1/CLK DFFPOSX1_46/D gnd vdd DFFPOSX1
XDFFPOSX1_24 BUFX2_26/A CLKBUF1_1/Y AOI22X1_54/Y gnd vdd DFFPOSX1
XAOI21X1_347 NOR2X1_36/Y BUFX4_152/Y BUFX4_14/Y gnd NAND2X1_622/A vdd AOI21X1
XAOI21X1_369 NAND2X1_571/Y NAND2X1_575/Y BUFX4_179/Y gnd OAI21X1_870/B vdd AOI21X1
XAOI21X1_336 OAI21X1_817/Y OAI21X1_813/Y OAI21X1_822/Y gnd AOI22X1_40/C vdd AOI21X1
XDFFPOSX1_13 BUFX2_15/A CLKBUF1_7/Y OAI21X1_843/Y gnd vdd DFFPOSX1
XAOI21X1_358 OR2X2_45/B BUFX4_60/Y NOR2X1_475/Y gnd NAND3X1_68/C vdd AOI21X1
XINVX1_162 INVX1_162/A gnd INVX1_162/Y vdd INVX1
XINVX1_184 operand_B[46] gnd INVX1_184/Y vdd INVX1
XINVX1_173 operand_B[43] gnd INVX1_173/Y vdd INVX1
XINVX1_140 INVX1_140/A gnd INVX1_140/Y vdd INVX1
XNAND2X1_509 BUFX4_70/Y OAI21X1_614/B gnd OAI21X1_592/C vdd NAND2X1
XINVX1_151 INVX1_151/A gnd INVX1_151/Y vdd INVX1
XINVX1_195 INVX1_195/A gnd OAI22X1_8/B vdd INVX1
XAOI21X1_111 INVX1_142/A NOR2X1_181/Y OAI21X1_357/Y gnd OAI21X1_358/C vdd AOI21X1
XAOI21X1_166 INVX1_199/Y OAI21X1_169/C OAI21X1_477/Y gnd OAI21X1_565/A vdd AOI21X1
XAOI21X1_133 OR2X2_21/B OR2X2_21/A BUFX4_94/Y gnd AOI21X1_136/A vdd AOI21X1
XFILL_20_2_0 gnd vdd FILL
XAOI21X1_100 OR2X2_7/B OAI21X1_333/Y AND2X2_14/Y gnd OR2X2_14/A vdd AOI21X1
XAOI21X1_144 BUFX4_163/Y MUX2X1_40/Y INVX8_15/Y gnd OAI21X1_435/C vdd AOI21X1
XAOI21X1_155 MUX2X1_34/S INVX1_54/A NOR2X1_235/Y gnd INVX1_189/A vdd AOI21X1
XAOI21X1_122 NOR2X1_75/A NOR2X1_197/Y AND2X2_18/Y gnd NOR2X1_198/B vdd AOI21X1
XAOI21X1_177 INVX4_23/Y NOR2X1_272/B BUFX4_32/Y gnd OAI21X1_498/C vdd AOI21X1
XAOI21X1_199 AND2X2_32/Y INVX1_223/Y INVX1_222/A gnd OAI21X1_563/A vdd AOI21X1
XAOI21X1_188 BUFX4_113/Y OAI22X1_30/D NAND3X1_30/Y gnd NAND2X1_459/A vdd AOI21X1
XFILL_28_3_0 gnd vdd FILL
XFILL_3_3_0 gnd vdd FILL
XFILL_11_2_0 gnd vdd FILL
XFILL_19_3_0 gnd vdd FILL
XBUFX4_9 BUFX4_9/A gnd BUFX4_9/Y vdd BUFX4
XNAND2X1_306 operand_A[36] operand_B[36] gnd INVX2_63/A vdd NAND2X1
XNAND2X1_317 MUX2X1_51/S OAI21X1_183/Y gnd OAI21X1_300/C vdd NAND2X1
XNAND2X1_339 MUX2X1_25/S MUX2X1_49/B gnd OAI21X1_326/C vdd NAND2X1
XNAND2X1_328 BUFX4_164/Y MUX2X1_34/B gnd OAI21X1_313/C vdd NAND2X1
XNOR2X1_394 NOR2X1_394/A NOR2X1_394/B gnd AND2X2_45/A vdd NOR2X1
XNOR2X1_383 BUFX2_45/A BUFX2_46/A gnd NOR2X1_383/Y vdd NOR2X1
XNOR2X1_350 NOR2X1_350/A BUFX4_145/Y gnd NOR2X1_351/A vdd NOR2X1
XNOR2X1_372 INVX4_18/A INVX1_74/Y gnd NOR2X1_372/Y vdd NOR2X1
XNOR2X1_361 BUFX4_163/Y NOR2X1_361/B gnd NOR2X1_361/Y vdd NOR2X1
XINVX4_9 operand_A[58] gnd INVX4_9/Y vdd INVX4
XOAI21X1_889 OAI21X1_889/A AOI22X1_50/Y AOI22X1_51/Y gnd NOR2X1_492/B vdd OAI21X1
XOAI21X1_867 NOR2X1_252/B NOR2X1_87/B OR2X2_40/B gnd OAI22X1_28/B vdd OAI21X1
XOAI21X1_834 INVX1_314/A NAND2X1_40/B BUFX4_140/Y gnd OAI21X1_834/Y vdd OAI21X1
XOAI21X1_845 INVX1_314/A NAND2X1_40/B NAND2X1_39/A gnd XNOR2X1_41/A vdd OAI21X1
XOAI21X1_823 XNOR2X1_6/Y OAI21X1_823/B OAI21X1_823/C gnd AOI22X1_42/D vdd OAI21X1
XOAI21X1_856 OAI21X1_856/A BUFX4_11/Y OAI21X1_856/C gnd OAI21X1_856/Y vdd OAI21X1
XOAI21X1_812 XNOR2X1_7/Y INVX2_93/Y OAI21X1_812/C gnd AOI22X1_40/D vdd OAI21X1
XOAI21X1_801 INVX8_15/Y OR2X2_43/Y OAI21X1_801/C gnd NOR2X1_453/B vdd OAI21X1
XOAI21X1_878 BUFX4_155/Y XNOR2X1_14/Y BUFX4_100/Y gnd NOR2X1_488/A vdd OAI21X1
XNOR2X1_90 INVX1_27/Y INVX2_36/Y gnd BUFX4_60/A vdd NOR2X1
XOAI21X1_119 INVX2_15/Y MUX2X1_6/S OAI21X1_119/C gnd INVX1_102/A vdd OAI21X1
XOAI21X1_108 INVX1_62/Y BUFX4_119/Y OAI21X1_108/C gnd INVX1_64/A vdd OAI21X1
XNAND2X1_114 BUFX4_50/Y operand_A[55] gnd OAI21X1_63/C vdd NAND2X1
XNAND2X1_125 BUFX4_184/Y OAI21X1_74/Y gnd OAI21X1_86/C vdd NAND2X1
XBUFX2_6 BUFX2_6/A gnd result[3] vdd BUFX2
XNAND2X1_103 BUFX4_74/Y INVX1_44/Y gnd OAI21X1_54/C vdd NAND2X1
XNAND2X1_1 operand_A[29] INVX2_1/Y gnd NAND2X1_3/A vdd NAND2X1
XNAND2X1_147 MUX2X1_4/S operand_A[24] gnd OAI21X1_102/C vdd NAND2X1
XNAND2X1_169 MUX2X1_99/S OAI21X1_272/A gnd OAI21X1_128/C vdd NAND2X1
XNAND2X1_136 OR2X2_13/B OAI21X1_84/Y gnd OAI21X1_85/C vdd NAND2X1
XNAND2X1_158 INVX8_1/A OAI21X1_113/Y gnd OAI21X1_114/C vdd NAND2X1
XNOR2X1_180 NOR2X1_185/A INVX1_156/A gnd INVX1_154/A vdd NOR2X1
XNOR2X1_191 INVX1_154/A INVX1_162/A gnd AND2X2_17/B vdd NOR2X1
XFILL_25_1_0 gnd vdd FILL
XFILL_0_1_0 gnd vdd FILL
XINVX2_6 operand_A[16] gnd INVX2_6/Y vdd INVX2
XOAI21X1_664 INVX2_65/Y OAI21X1_664/B OAI21X1_664/C gnd NOR2X1_421/A vdd OAI21X1
XOAI21X1_620 OAI22X1_22/D INVX2_91/A OAI21X1_626/A gnd NAND3X1_37/C vdd OAI21X1
XOAI21X1_653 NOR2X1_67/A NAND2X1_50/B AOI22X1_1/A gnd OAI21X1_653/Y vdd OAI21X1
XOAI21X1_675 OAI21X1_675/A NOR2X1_413/Y OAI21X1_675/C gnd AOI22X1_31/C vdd OAI21X1
XMUX2X1_120 MUX2X1_120/A MUX2X1_120/B BUFX4_16/Y gnd NOR2X1_458/B vdd MUX2X1
XOAI21X1_631 OAI21X1_631/A BUFX4_25/Y MUX2X1_49/S gnd OAI22X1_23/B vdd OAI21X1
XOAI21X1_642 INVX2_58/Y INVX1_279/Y AOI21X1_48/A gnd OAI21X1_643/A vdd OAI21X1
XOAI21X1_686 INVX2_16/Y MUX2X1_4/S OAI21X1_36/C gnd OAI21X1_686/Y vdd OAI21X1
XAOI21X1_6 INVX2_10/Y XOR2X1_3/Y NOR2X1_15/Y gnd OAI21X1_9/A vdd AOI21X1
XOAI21X1_697 OAI22X1_7/C NOR2X1_409/A BUFX4_97/Y gnd OAI21X1_697/Y vdd OAI21X1
XXNOR2X1_36 XNOR2X1_36/A INVX1_204/A gnd XNOR2X1_36/Y vdd XNOR2X1
XXNOR2X1_47 XNOR2X1_47/A XNOR2X1_47/B gnd XNOR2X1_47/Y vdd XNOR2X1
XINVX1_60 INVX1_60/A gnd INVX1_60/Y vdd INVX1
XFILL_8_2_0 gnd vdd FILL
XXNOR2X1_25 operand_B[16] operand_A[16] gnd XNOR2X1_25/Y vdd XNOR2X1
XXNOR2X1_14 operand_A[18] operand_B[18] gnd XNOR2X1_14/Y vdd XNOR2X1
XBUFX2_46 BUFX2_46/A gnd result[43] vdd BUFX2
XBUFX2_57 OR2X2_37/A gnd result[54] vdd BUFX2
XBUFX2_35 BUFX2_35/A gnd result[32] vdd BUFX2
XINVX1_71 INVX1_71/A gnd INVX1_71/Y vdd INVX1
XFILL_16_1_0 gnd vdd FILL
XDFFPOSX1_1 BUFX2_3/A DFFSR_1/CLK DFFPOSX1_1/D gnd vdd DFFPOSX1
XBUFX2_24 OR2X2_48/B gnd result[21] vdd BUFX2
XINVX1_82 INVX1_82/A gnd INVX1_82/Y vdd INVX1
XBUFX2_13 BUFX2_13/A gnd result[10] vdd BUFX2
XINVX1_93 INVX1_93/A gnd INVX1_93/Y vdd INVX1
XNOR2X1_4 operand_B[22] INVX4_3/Y gnd NOR2X1_4/Y vdd NOR2X1
XAOI21X1_69 NAND3X1_6/Y AOI21X1_69/B NOR2X1_133/Y gnd AOI21X1_69/Y vdd AOI21X1
XAOI21X1_47 NOR2X1_106/Y INVX1_315/A AOI21X1_47/C gnd INVX1_77/A vdd AOI21X1
XAOI21X1_36 BUFX4_81/Y OAI21X1_86/Y INVX8_9/Y gnd OAI22X1_2/C vdd AOI21X1
XAOI21X1_58 NOR2X1_48/Y OAI21X1_26/Y INVX1_28/A gnd AOI21X1_58/Y vdd AOI21X1
XAOI21X1_25 NOR2X1_58/Y XNOR2X1_18/Y INVX1_81/A gnd OAI21X1_29/C vdd AOI21X1
XAOI21X1_14 OAI21X1_17/Y NOR2X1_29/Y OAI21X1_18/Y gnd OAI21X1_19/C vdd AOI21X1
XOAI21X1_9 OAI21X1_9/A OAI21X1_9/B OAI21X1_9/C gnd OAI21X1_9/Y vdd OAI21X1
XOAI22X1_11 BUFX4_157/Y INVX2_78/Y BUFX4_145/Y OAI22X1_11/D gnd OAI22X1_11/Y vdd OAI22X1
XOAI22X1_22 BUFX4_64/Y INVX2_91/Y BUFX4_145/Y OAI22X1_22/D gnd OAI22X1_22/Y vdd OAI22X1
XOAI21X1_450 operand_A[45] operand_B[45] AND2X2_21/Y gnd OAI21X1_451/C vdd OAI21X1
XOAI22X1_33 BUFX4_81/Y OAI22X1_33/B OAI22X1_33/C OAI22X1_33/D gnd OAI22X1_33/Y vdd
+ OAI22X1
XOAI21X1_472 INVX1_77/A OAI21X1_472/B OAI21X1_472/C gnd AND2X2_26/A vdd OAI21X1
XOAI21X1_461 OAI22X1_7/C NOR2X1_231/A AOI22X1_16/Y gnd OR2X2_26/A vdd OAI21X1
XOAI21X1_483 INVX8_7/Y MUX2X1_42/Y NOR2X1_253/Y gnd OAI21X1_483/Y vdd OAI21X1
XOAI21X1_494 OAI22X1_1/B NAND3X1_7/Y OAI21X1_494/C gnd OAI21X1_494/Y vdd OAI21X1
XFILL_32_4_1 gnd vdd FILL
XFILL_23_4_1 gnd vdd FILL
XBUFX4_108 NOR2X1_45/Y gnd BUFX4_108/Y vdd BUFX4
XFILL_5_0_0 gnd vdd FILL
XBUFX4_119 INVX8_3/Y gnd BUFX4_119/Y vdd BUFX4
XFILL_6_5_1 gnd vdd FILL
XFILL_14_4_1 gnd vdd FILL
XOAI21X1_280 INVX1_59/Y BUFX4_133/Y OAI21X1_280/C gnd OAI21X1_411/B vdd OAI21X1
XOAI21X1_291 MUX2X1_87/S INVX1_92/A OAI21X1_291/C gnd MUX2X1_31/A vdd OAI21X1
XINVX1_300 OR2X2_40/Y gnd INVX1_300/Y vdd INVX1
XINVX1_322 BUFX2_28/A gnd INVX1_322/Y vdd INVX1
XINVX1_311 NOR2X1_37/Y gnd INVX1_311/Y vdd INVX1
XFILL_29_1 gnd vdd FILL
XAOI21X1_315 BUFX4_81/Y MUX2X1_107/Y INVX8_9/Y gnd OAI22X1_27/B vdd AOI21X1
XAOI21X1_304 XOR2X1_3/Y NOR2X1_112/Y BUFX4_92/Y gnd OAI21X1_713/C vdd AOI21X1
XAOI21X1_326 XOR2X1_5/Y OAI21X1_782/B BUFX4_27/Y gnd OAI21X1_782/C vdd AOI21X1
XAOI21X1_337 XOR2X1_8/Y INVX2_93/A NOR2X1_35/Y gnd OAI21X1_823/B vdd AOI21X1
XAOI21X1_348 BUFX4_85/Y NOR2X1_227/Y NAND2X1_622/Y gnd NAND3X1_66/A vdd AOI21X1
XDFFPOSX1_58 OR2X2_37/B CLKBUF1_5/Y DFFPOSX1_58/D gnd vdd DFFPOSX1
XDFFPOSX1_36 BUFX2_38/A CLKBUF1_3/Y AOI21X1_81/Y gnd vdd DFFPOSX1
XDFFPOSX1_47 BUFX2_49/A CLKBUF1_8/Y DFFPOSX1_47/D gnd vdd DFFPOSX1
XDFFPOSX1_25 BUFX2_27/A CLKBUF1_1/Y DFFPOSX1_25/D gnd vdd DFFPOSX1
XAOI21X1_359 INVX1_313/Y AOI21X1_359/B NAND3X1_68/Y gnd OAI21X1_856/A vdd AOI21X1
XDFFPOSX1_14 BUFX2_16/A CLKBUF1_7/Y DFFPOSX1_14/D gnd vdd DFFPOSX1
XINVX1_141 OR2X2_36/A gnd INVX1_141/Y vdd INVX1
XINVX1_152 operand_B[40] gnd INVX1_152/Y vdd INVX1
XINVX1_130 INVX1_130/A gnd INVX1_130/Y vdd INVX1
XINVX1_163 INVX1_163/A gnd INVX1_163/Y vdd INVX1
XINVX1_185 INVX1_185/A gnd OR2X2_28/B vdd INVX1
XINVX1_174 INVX1_174/A gnd INVX1_174/Y vdd INVX1
XINVX1_196 INVX1_196/A gnd INVX1_196/Y vdd INVX1
XNOR2X1_510 NOR2X1_510/A NOR2X1_510/B gnd NOR2X1_510/Y vdd NOR2X1
XAOI21X1_167 AND2X2_26/B OAI21X1_565/A BUFX4_93/Y gnd OAI21X1_478/C vdd AOI21X1
XAOI21X1_189 BUFX4_143/Y XNOR2X1_38/Y NAND2X1_459/Y gnd AOI21X1_190/A vdd AOI21X1
XAOI21X1_123 OAI21X1_380/Y NOR2X1_192/Y NAND3X1_18/Y gnd AOI21X1_124/B vdd AOI21X1
XAOI21X1_112 INVX1_154/Y INVX1_155/Y BUFX4_28/Y gnd AOI21X1_115/B vdd AOI21X1
XAOI21X1_178 INVX1_200/A OAI21X1_362/Y OAI21X1_499/Y gnd OAI21X1_500/C vdd AOI21X1
XAOI21X1_134 INVX8_17/A NOR2X1_210/B OAI22X1_7/Y gnd NAND2X1_394/B vdd AOI21X1
XAOI21X1_145 OAI21X1_425/Y NOR2X1_221/Y OR2X2_23/Y gnd AOI21X1_146/B vdd AOI21X1
XFILL_20_2_1 gnd vdd FILL
XAOI21X1_156 INVX4_20/A INVX1_189/Y OR2X2_26/Y gnd NAND3X1_25/C vdd AOI21X1
XAOI21X1_101 NOR2X1_75/A OAI21X1_342/Y AND2X2_14/Y gnd OAI21X1_780/A vdd AOI21X1
XFILL_28_3_1 gnd vdd FILL
XFILL_3_3_1 gnd vdd FILL
XFILL_11_2_1 gnd vdd FILL
XFILL_19_3_1 gnd vdd FILL
XNAND2X1_307 operand_B[35] INVX2_61/Y gnd AOI21X1_84/A vdd NAND2X1
XNAND2X1_318 BUFX4_159/Y MUX2X1_33/Y gnd OAI21X1_304/C vdd NAND2X1
XNAND2X1_329 BUFX4_122/Y OAI21X1_231/B gnd OAI21X1_311/C vdd NAND2X1
XNOR2X1_384 OR2X2_36/Y NOR2X1_384/B gnd NOR2X1_384/Y vdd NOR2X1
XNOR2X1_340 operand_B[58] INVX4_9/Y gnd NOR2X1_341/A vdd NOR2X1
XNOR2X1_351 NOR2X1_351/A OAI22X1_20/Y gnd AND2X2_43/A vdd NOR2X1
XNOR2X1_362 OR2X2_8/B NOR2X1_362/B gnd NOR2X1_362/Y vdd NOR2X1
XNOR2X1_373 BUFX4_36/Y NOR2X1_373/B gnd OAI22X1_23/A vdd NOR2X1
XNOR2X1_395 BUFX2_16/A BUFX2_15/A gnd NOR2X1_395/Y vdd NOR2X1
XOAI21X1_813 OR2X2_19/A BUFX4_9/Y OAI21X1_813/C gnd OAI21X1_813/Y vdd OAI21X1
XOAI21X1_835 OAI21X1_835/A INVX1_309/Y OAI21X1_835/C gnd OAI21X1_842/B vdd OAI21X1
XOAI21X1_824 operand_B[10] INVX2_22/Y OAI21X1_824/C gnd OAI21X1_825/B vdd OAI21X1
XOAI21X1_857 XNOR2X1_22/Y NOR2X1_476/Y OAI21X1_857/C gnd OAI21X1_857/Y vdd OAI21X1
XOAI21X1_846 NOR2X1_470/Y NOR2X1_471/Y MUX2X1_64/S gnd OAI21X1_848/C vdd OAI21X1
XOAI21X1_802 OAI21X1_802/A OR2X2_42/Y BUFX4_100/Y gnd OAI21X1_803/C vdd OAI21X1
XOAI21X1_868 INVX4_26/Y OR2X2_46/Y OAI21X1_868/C gnd AOI22X1_47/D vdd OAI21X1
XOAI21X1_879 INVX4_5/Y INVX2_5/Y NAND3X1_70/B gnd OAI21X1_880/B vdd OAI21X1
XNOR2X1_91 NOR2X1_91/A NOR2X1_91/B gnd NOR2X1_91/Y vdd NOR2X1
XNOR2X1_80 NOR2X1_80/A INVX4_10/Y gnd INVX4_11/A vdd NOR2X1
XBUFX2_7 BUFX2_7/A gnd result[4] vdd BUFX2
XOAI21X1_109 BUFX4_23/Y OAI21X1_109/B OAI21X1_109/C gnd AND2X2_25/A vdd OAI21X1
XFILL_11_1 gnd vdd FILL
XNAND2X1_137 operand_A[31] operand_B[31] gnd INVX1_75/A vdd NAND2X1
XNAND2X1_126 MUX2X1_1/S operand_A[37] gnd OAI21X1_75/C vdd NAND2X1
XNAND2X1_115 MUX2X1_7/S operand_A[57] gnd OAI21X1_64/C vdd NAND2X1
XNAND2X1_148 BUFX4_46/Y operand_A[26] gnd OAI21X1_704/C vdd NAND2X1
XNAND2X1_104 MUX2X1_8/S operand_A[11] gnd OAI21X1_55/C vdd NAND2X1
XNAND2X1_159 BUFX4_125/Y INVX1_122/A gnd OAI21X1_115/C vdd NAND2X1
XNAND2X1_2 operand_B[29] INVX2_2/Y gnd AND2X2_2/B vdd NAND2X1
XFILL_25_1_1 gnd vdd FILL
XNOR2X1_181 OR2X2_12/B INVX1_148/A gnd NOR2X1_181/Y vdd NOR2X1
XNOR2X1_192 NOR2X1_192/A AND2X2_17/Y gnd NOR2X1_192/Y vdd NOR2X1
XOAI21X1_621 OAI21X1_621/A OAI21X1_621/B INVX1_259/A gnd NAND3X1_38/C vdd OAI21X1
XOAI21X1_610 OAI21X1_610/A INVX1_248/A INVX1_253/Y gnd OAI21X1_610/Y vdd OAI21X1
XOAI21X1_632 INVX8_7/Y OAI22X1_23/Y NOR2X1_372/Y gnd OAI21X1_633/C vdd OAI21X1
XFILL_0_1_1 gnd vdd FILL
XNOR2X1_170 INVX8_8/Y NOR2X1_170/B gnd OAI22X1_6/B vdd NOR2X1
XINVX2_7 operand_A[19] gnd INVX2_7/Y vdd INVX2
XOAI21X1_665 INVX2_62/Y OAI21X1_665/B AOI21X1_84/A gnd OAI21X1_665/Y vdd OAI21X1
XOAI21X1_654 OAI21X1_654/A NOR2X1_121/B OAI21X1_654/C gnd OAI21X1_654/Y vdd OAI21X1
XOAI21X1_676 INVX2_31/Y MUX2X1_5/S OAI21X1_46/C gnd OAI21X1_676/Y vdd OAI21X1
XMUX2X1_121 MUX2X1_33/B MUX2X1_121/B BUFX4_39/Y gnd MUX2X1_129/B vdd MUX2X1
XOAI21X1_643 OAI21X1_643/A OAI21X1_28/A OAI21X1_643/C gnd AND2X2_47/A vdd OAI21X1
XOAI21X1_687 INVX1_288/Y NOR2X1_54/A OAI21X1_687/C gnd MUX2X1_106/A vdd OAI21X1
XMUX2X1_110 MUX2X1_110/A MUX2X1_110/B NOR2X1_19/B gnd MUX2X1_110/Y vdd MUX2X1
XAOI21X1_7 NOR2X1_17/Y XOR2X1_4/Y NOR2X1_16/Y gnd OAI21X1_9/C vdd AOI21X1
XOAI21X1_698 INVX1_100/A INVX8_15/Y AND2X2_51/Y gnd OAI21X1_698/Y vdd OAI21X1
XXNOR2X1_37 XNOR2X1_37/A INVX4_23/Y gnd XNOR2X1_37/Y vdd XNOR2X1
XXNOR2X1_48 XNOR2X1_48/A NOR2X1_67/A gnd XNOR2X1_48/Y vdd XNOR2X1
XXNOR2X1_26 operand_B[27] operand_A[27] gnd XNOR2X1_26/Y vdd XNOR2X1
XINVX1_72 INVX1_72/A gnd INVX1_72/Y vdd INVX1
XINVX1_50 INVX1_50/A gnd INVX1_50/Y vdd INVX1
XINVX1_61 INVX1_61/A gnd INVX1_61/Y vdd INVX1
XINVX1_83 INVX1_83/A gnd INVX1_83/Y vdd INVX1
XFILL_8_2_1 gnd vdd FILL
XXNOR2X1_15 operand_B[19] operand_A[19] gnd XNOR2X1_15/Y vdd XNOR2X1
XINVX1_94 INVX1_94/A gnd INVX1_94/Y vdd INVX1
XBUFX2_36 BUFX2_36/A gnd result[33] vdd BUFX2
XBUFX2_58 BUFX2_58/A gnd result[55] vdd BUFX2
XBUFX2_47 BUFX2_47/A gnd result[44] vdd BUFX2
XBUFX2_25 BUFX2_25/A gnd result[22] vdd BUFX2
XFILL_16_1_1 gnd vdd FILL
XBUFX2_14 BUFX2_14/A gnd result[11] vdd BUFX2
XDFFPOSX1_2 BUFX2_4/A DFFSR_1/CLK DFFPOSX1_2/D gnd vdd DFFPOSX1
XNOR2X1_5 operand_B[21] INVX4_4/Y gnd NOR2X1_5/Y vdd NOR2X1
XAOI21X1_37 OAI21X1_24/Y NOR2X1_91/Y NOR2X1_92/Y gnd AOI21X1_37/Y vdd AOI21X1
XAOI21X1_59 NOR2X1_97/A OAI21X1_94/C NOR2X1_123/Y gnd AOI21X1_59/Y vdd AOI21X1
XAOI21X1_15 AND2X2_1/Y INVX1_315/A INVX1_10/Y gnd OAI21X1_23/A vdd AOI21X1
XAOI21X1_48 AOI21X1_48/A INVX1_279/A INVX2_10/A gnd NOR2X1_428/A vdd AOI21X1
XAOI21X1_26 NOR2X1_56/Y OAI21X1_28/Y OAI21X1_29/Y gnd OAI21X1_32/A vdd AOI21X1
XOAI22X1_12 OR2X2_16/B OAI22X1_12/B MUX2X1_48/Y INVX8_7/Y gnd OAI22X1_12/Y vdd OAI22X1
XOAI22X1_34 OAI22X1_34/A OAI22X1_34/B OAI22X1_34/C OAI22X1_34/D gnd OAI22X1_34/Y vdd
+ OAI22X1
XOAI22X1_23 OAI22X1_23/A OAI22X1_23/B OAI22X1_23/C MUX2X1_49/S gnd OAI22X1_23/Y vdd
+ OAI22X1
XOAI21X1_473 AND2X2_26/B AND2X2_26/A NOR2X1_246/Y gnd OAI21X1_473/Y vdd OAI21X1
XOAI21X1_462 NOR2X1_231/B NOR2X1_231/A OR2X2_24/A gnd NAND3X1_26/C vdd OAI21X1
XOAI21X1_451 INVX4_14/Y INVX1_179/Y OAI21X1_451/C gnd INVX1_185/A vdd OAI21X1
XOAI21X1_440 INVX4_14/Y MUX2X1_5/S OAI21X1_440/C gnd INVX1_180/A vdd OAI21X1
XOAI21X1_484 INVX1_99/Y BUFX4_41/Y BUFX4_186/Y gnd OAI21X1_485/C vdd OAI21X1
XOAI21X1_495 operand_A[49] operand_B[49] BUFX4_4/Y gnd AND2X2_29/B vdd OAI21X1
XNAND2X1_490 NOR2X1_310/Y OAI21X1_546/Y gnd NAND2X1_492/B vdd NAND2X1
XBUFX4_109 operand_B[5] gnd NOR2X1_22/A vdd BUFX4
XFILL_5_0_1 gnd vdd FILL
XOAI21X1_270 BUFX4_63/Y OAI21X1_283/C AOI22X1_6/Y gnd NOR2X1_148/B vdd OAI21X1
XINVX1_323 NOR2X1_42/Y gnd INVX1_323/Y vdd INVX1
XINVX1_312 INVX1_312/A gnd INVX1_312/Y vdd INVX1
XINVX1_301 INVX1_301/A gnd INVX1_301/Y vdd INVX1
XOAI21X1_281 INVX1_123/Y BUFX4_20/Y OAI21X1_281/C gnd INVX1_124/A vdd OAI21X1
XOAI21X1_292 INVX1_128/Y BUFX4_119/Y OAI21X1_292/C gnd INVX1_129/A vdd OAI21X1
XAND2X2_70 AND2X2_70/A AND2X2_70/B gnd AND2X2_70/Y vdd AND2X2
XAOI21X1_316 XNOR2X1_21/Y OAI21X1_28/Y BUFX4_92/Y gnd OAI21X1_752/C vdd AOI21X1
XAOI21X1_338 XNOR2X1_6/Y OAI21X1_823/B BUFX4_31/Y gnd OAI21X1_823/C vdd AOI21X1
XAOI21X1_327 AOI21X1_9/Y INVX1_17/A OAI21X1_793/Y gnd OR2X2_42/B vdd AOI21X1
XAOI21X1_305 BUFX4_162/Y MUX2X1_96/Y OAI21X1_728/Y gnd NOR2X1_433/B vdd AOI21X1
XAOI21X1_349 BUFX4_140/Y XNOR2X1_41/Y NAND3X1_66/Y gnd AOI21X1_350/B vdd AOI21X1
XDFFPOSX1_37 BUFX2_39/A CLKBUF1_3/Y OAI21X1_306/Y gnd vdd DFFPOSX1
XDFFPOSX1_59 BUFX2_61/A CLKBUF1_5/Y DFFPOSX1_59/D gnd vdd DFFPOSX1
XDFFPOSX1_48 BUFX2_50/A CLKBUF1_8/Y DFFPOSX1_48/D gnd vdd DFFPOSX1
XDFFPOSX1_26 BUFX2_28/A CLKBUF1_1/Y OAI21X1_920/Y gnd vdd DFFPOSX1
XDFFPOSX1_15 BUFX2_17/A CLKBUF1_2/Y OAI21X1_856/Y gnd vdd DFFPOSX1
XINVX1_142 INVX1_142/A gnd INVX1_142/Y vdd INVX1
XINVX1_153 INVX1_153/A gnd INVX1_153/Y vdd INVX1
XINVX1_186 INVX1_186/A gnd OR2X2_24/B vdd INVX1
XINVX1_164 INVX1_164/A gnd INVX1_164/Y vdd INVX1
XINVX1_131 INVX1_131/A gnd INVX1_131/Y vdd INVX1
XINVX1_175 INVX1_175/A gnd INVX1_175/Y vdd INVX1
XINVX1_120 INVX1_120/A gnd INVX1_120/Y vdd INVX1
XINVX1_197 operand_B[48] gnd INVX1_197/Y vdd INVX1
XNOR2X1_511 NOR2X1_93/A BUFX2_32/A gnd NOR2X1_511/Y vdd NOR2X1
XNOR2X1_500 NOR2X1_500/A NOR2X1_500/B gnd NOR2X1_500/Y vdd NOR2X1
XAOI21X1_102 INVX1_148/Y OAI21X1_347/B BUFX4_28/Y gnd OAI21X1_347/C vdd AOI21X1
XAOI21X1_124 OAI21X1_379/Y AOI21X1_124/B NOR2X1_187/Y gnd DFFPOSX1_42/D vdd AOI21X1
XAOI21X1_179 NOR2X1_265/Y OAI21X1_500/Y OAI21X1_501/Y gnd XNOR2X1_37/A vdd AOI21X1
XAOI21X1_146 OAI21X1_423/Y AOI21X1_146/B NOR2X1_215/Y gnd DFFPOSX1_45/D vdd AOI21X1
XAOI21X1_113 INVX1_158/Y OAI21X1_169/C OAI21X1_362/Y gnd INVX1_163/A vdd AOI21X1
XAOI21X1_157 OR2X2_24/Y NOR2X1_234/Y NAND3X1_25/Y gnd AOI21X1_158/B vdd AOI21X1
XAOI21X1_168 INVX4_11/Y NOR2X1_252/B BUFX4_7/Y gnd OAI22X1_28/A vdd AOI21X1
XAOI21X1_135 INVX4_18/A NOR2X1_213/Y NAND2X1_394/Y gnd NAND3X1_20/A vdd AOI21X1
XFILL_30_5_0 gnd vdd FILL
XNAND2X1_319 MUX2X1_30/S OAI21X1_177/B gnd OAI21X1_301/C vdd NAND2X1
XNAND2X1_308 MUX2X1_2/S OAI21X1_187/Y gnd OAI21X1_290/C vdd NAND2X1
XNOR2X1_385 BUFX2_55/A BUFX2_56/A gnd NOR2X1_385/Y vdd NOR2X1
XNOR2X1_363 BUFX4_98/Y BUFX2_64/A gnd NOR2X1_363/Y vdd NOR2X1
XNOR2X1_341 NOR2X1_341/A AND2X2_41/Y gnd NOR2X1_341/Y vdd NOR2X1
XNOR2X1_330 INVX2_81/Y INVX2_82/Y gnd INVX1_239/A vdd NOR2X1
XNOR2X1_374 NOR2X1_374/A NOR2X1_374/B gnd NOR2X1_374/Y vdd NOR2X1
XNOR2X1_352 NOR2X1_352/A NOR2X1_352/B gnd NOR2X1_352/Y vdd NOR2X1
XFILL_21_5_0 gnd vdd FILL
XOAI21X1_814 BUFX4_35/Y MUX2X1_96/A OAI21X1_814/C gnd OAI21X1_815/A vdd OAI21X1
XNOR2X1_396 BUFX2_10/A BUFX2_9/A gnd NOR2X1_396/Y vdd NOR2X1
XOAI21X1_803 OR2X2_48/A INVX1_265/Y OAI21X1_803/C gnd DFFPOSX1_9/D vdd OAI21X1
XOAI21X1_858 OR2X2_45/A INVX2_19/Y INVX2_18/A gnd OAI21X1_859/A vdd OAI21X1
XOAI21X1_825 XNOR2X1_6/Y OAI21X1_825/B OAI21X1_825/C gnd AND2X2_60/B vdd OAI21X1
XOAI21X1_869 NOR2X1_485/B OAI21X1_7/C NAND2X1_19/A gnd XNOR2X1_42/A vdd OAI21X1
XOAI21X1_847 OAI21X1_847/A BUFX4_24/Y OAI21X1_847/C gnd INVX1_328/A vdd OAI21X1
XOAI21X1_836 NOR2X1_465/Y NOR2X1_464/Y MUX2X1_25/S gnd AND2X2_61/A vdd OAI21X1
XFILL_12_5_0 gnd vdd FILL
XNAND3X1_70 BUFX4_108/Y NAND3X1_70/B OR2X2_47/Y gnd NAND3X1_70/Y vdd NAND3X1
XNOR2X1_92 BUFX2_33/A NOR2X1_93/A gnd NOR2X1_92/Y vdd NOR2X1
XNOR2X1_70 NOR2X1_70/A NOR2X1_70/B gnd INVX1_33/A vdd NOR2X1
XNOR2X1_81 INVX4_10/Y BUFX4_21/Y gnd INVX2_48/A vdd NOR2X1
XBUFX2_8 BUFX2_8/A gnd result[5] vdd BUFX2
XNAND2X1_138 INVX2_50/Y INVX2_51/Y gnd AND2X2_6/A vdd NAND2X1
XNAND2X1_3 NAND2X1_3/A AND2X2_2/B gnd NAND2X1_3/Y vdd NAND2X1
XNAND2X1_127 BUFX4_71/Y MUX2X1_6/Y gnd OAI21X1_76/C vdd NAND2X1
XNAND2X1_116 INVX8_1/A MUX2X1_22/A gnd OAI21X1_65/C vdd NAND2X1
XNAND2X1_149 BUFX4_69/Y OAI21X1_103/Y gnd OAI21X1_104/C vdd NAND2X1
XNAND2X1_105 BUFX4_191/Y OAI21X1_55/Y gnd OAI21X1_56/C vdd NAND2X1
XNOR2X1_160 INVX8_8/Y INVX1_132/Y gnd OAI22X1_27/A vdd NOR2X1
XOAI21X1_600 INVX2_88/A OAI21X1_600/B NOR2X1_347/Y gnd OAI21X1_600/Y vdd OAI21X1
XNOR2X1_182 NOR2X1_420/A NOR2X1_183/B gnd INVX1_157/A vdd NOR2X1
XOAI21X1_611 INVX1_257/A INVX1_255/A INVX2_88/Y gnd OR2X2_38/A vdd OAI21X1
XOAI21X1_666 INVX4_16/Y OAI21X1_666/B OAI21X1_666/C gnd OAI21X1_666/Y vdd OAI21X1
XOAI21X1_622 INVX4_12/Y operand_B[61] OAI21X1_622/C gnd INVX1_260/A vdd OAI21X1
XNOR2X1_171 NOR2X1_171/A NOR2X1_171/B gnd NOR2X1_171/Y vdd NOR2X1
XOAI21X1_655 NAND3X1_54/Y OAI21X1_655/B NOR2X1_412/Y gnd OAI21X1_655/Y vdd OAI21X1
XINVX2_8 operand_A[23] gnd INVX2_8/Y vdd INVX2
XOAI21X1_633 BUFX4_80/Y AOI21X1_41/C OAI21X1_633/C gnd NAND3X1_41/C vdd OAI21X1
XNOR2X1_193 BUFX4_179/Y MUX2X1_37/Y gnd NOR2X1_193/Y vdd NOR2X1
XAOI21X1_8 NOR2X1_26/Y XOR2X1_5/Y NOR2X1_25/Y gnd AOI21X1_8/Y vdd AOI21X1
XOAI21X1_644 OAI21X1_644/A OR2X2_3/A OAI21X1_644/C gnd OAI21X1_645/B vdd OAI21X1
XOAI21X1_677 BUFX4_191/Y MUX2X1_70/Y OAI21X1_677/C gnd MUX2X1_71/A vdd OAI21X1
XMUX2X1_111 MUX2X1_111/A MUX2X1_111/B MUX2X1_71/S gnd MUX2X1_112/A vdd MUX2X1
XOAI21X1_699 AND2X2_52/Y AOI21X1_66/Y INVX8_4/A gnd AND2X2_53/A vdd OAI21X1
XMUX2X1_100 MUX2X1_93/B MUX2X1_90/A BUFX4_66/Y gnd MUX2X1_113/A vdd MUX2X1
XOAI21X1_688 INVX1_287/Y MUX2X1_99/S OAI21X1_688/C gnd OAI21X1_796/B vdd OAI21X1
XMUX2X1_122 MUX2X1_122/A MUX2X1_122/B INVX8_2/A gnd MUX2X1_122/Y vdd MUX2X1
XXNOR2X1_38 XNOR2X1_38/A INVX1_212/A gnd XNOR2X1_38/Y vdd XNOR2X1
XXNOR2X1_49 XNOR2X1_49/A NAND2X1_3/Y gnd XNOR2X1_49/Y vdd XNOR2X1
XNAND2X1_650 NOR2X1_505/Y OAI22X1_38/Y gnd NOR2X1_506/B vdd NAND2X1
XXNOR2X1_27 operand_B[26] operand_A[26] gnd XNOR2X1_27/Y vdd XNOR2X1
XBUFX2_26 BUFX2_26/A gnd result[23] vdd BUFX2
XINVX1_95 INVX1_95/A gnd INVX1_95/Y vdd INVX1
XINVX1_51 INVX1_51/A gnd INVX1_51/Y vdd INVX1
XINVX1_73 INVX1_73/A gnd INVX1_73/Y vdd INVX1
XINVX1_84 INVX1_84/A gnd INVX1_84/Y vdd INVX1
XXNOR2X1_16 MUX2X1_99/S operand_A[2] gnd XNOR2X1_16/Y vdd XNOR2X1
XBUFX2_15 BUFX2_15/A gnd result[12] vdd BUFX2
XINVX1_62 INVX1_62/A gnd INVX1_62/Y vdd INVX1
XINVX1_40 INVX1_40/A gnd INVX1_40/Y vdd INVX1
XBUFX2_37 BUFX2_37/A gnd result[34] vdd BUFX2
XBUFX2_48 BUFX2_48/A gnd result[45] vdd BUFX2
XBUFX2_59 BUFX2_59/A gnd result[56] vdd BUFX2
XDFFPOSX1_3 BUFX2_5/A CLKBUF1_7/Y DFFPOSX1_3/D gnd vdd DFFPOSX1
XNOR2X1_6 NOR2X1_6/A NOR2X1_6/B gnd NOR2X1_6/Y vdd NOR2X1
XAOI21X1_16 NAND2X1_52/Y NOR2X1_42/Y NOR2X1_41/Y gnd OAI21X1_22/B vdd AOI21X1
XAOI21X1_38 OAI21X1_94/C NOR2X1_94/Y BUFX4_29/Y gnd OAI21X1_93/C vdd AOI21X1
XAOI21X1_49 OAI21X1_9/C AOI21X1_49/B NAND3X1_4/Y gnd AOI21X1_49/Y vdd AOI21X1
XAOI21X1_27 NAND2X1_79/Y NOR2X1_62/Y NOR2X1_61/Y gnd OAI21X1_30/B vdd AOI21X1
XOAI22X1_13 BUFX4_157/Y INVX1_224/Y BUFX4_145/Y OAI22X1_13/D gnd OAI22X1_13/Y vdd
+ OAI22X1
XFILL_26_4_0 gnd vdd FILL
XOAI22X1_24 INVX1_245/Y operand_A[60] operand_A[61] INVX1_252/Y gnd OAI22X1_24/Y vdd
+ OAI22X1
XOAI22X1_35 OAI22X1_35/A OAI22X1_35/B OAI22X1_35/C OAI22X1_35/D gnd OAI22X1_35/Y vdd
+ OAI22X1
XFILL_1_4_0 gnd vdd FILL
XOAI21X1_463 AND2X2_24/Y INVX1_192/A INVX4_22/A gnd NAND3X1_27/C vdd OAI21X1
XOAI21X1_452 NOR2X1_220/B NOR2X1_244/A OR2X2_28/B gnd OAI21X1_453/B vdd OAI21X1
XOAI21X1_430 OAI22X1_3/C NOR2X1_217/A AOI22X1_13/Y gnd NOR2X1_224/B vdd OAI21X1
XOAI21X1_474 NOR2X1_217/A AND2X2_21/Y INVX4_21/A gnd OR2X2_29/A vdd OAI21X1
XOAI21X1_441 INVX1_180/Y BUFX4_192/Y OAI21X1_441/C gnd OAI21X1_441/Y vdd OAI21X1
XOAI21X1_496 OAI21X1_871/A BUFX4_173/Y AND2X2_30/Y gnd OAI21X1_496/Y vdd OAI21X1
XOAI21X1_485 MUX2X1_25/B INVX8_5/A OAI21X1_485/C gnd NOR2X1_484/B vdd OAI21X1
XFILL_9_5_0 gnd vdd FILL
XNAND2X1_491 operand_B[55] INVX2_80/Y gnd OAI21X1_660/C vdd NAND2X1
XFILL_17_4_0 gnd vdd FILL
XNAND2X1_480 BUFX4_167/Y OAI21X1_342/Y gnd OAI21X1_903/A vdd NAND2X1
XOAI21X1_90 INVX1_54/Y BUFX4_186/Y INVX4_11/Y gnd AND2X2_3/A vdd OAI21X1
XOAI21X1_293 INVX2_44/Y BUFX4_46/Y OAI21X1_293/C gnd INVX1_130/A vdd OAI21X1
XINVX1_324 INVX1_324/A gnd INVX1_324/Y vdd INVX1
XOAI21X1_271 OR2X2_10/Y OR2X2_32/B NOR2X1_148/Y gnd NOR2X1_149/A vdd OAI21X1
XINVX1_302 INVX1_302/A gnd INVX1_302/Y vdd INVX1
XINVX1_313 INVX1_313/A gnd INVX1_313/Y vdd INVX1
XOAI21X1_282 INVX1_124/Y MUX2X1_25/S OAI21X1_282/C gnd AOI22X1_7/B vdd OAI21X1
XOAI21X1_260 INVX1_114/Y BUFX4_17/Y OAI21X1_260/C gnd OAI21X1_506/A vdd OAI21X1
XAND2X2_71 AND2X2_71/A AND2X2_71/B gnd AND2X2_71/Y vdd AND2X2
XAND2X2_60 AND2X2_60/A AND2X2_60/B gnd AND2X2_60/Y vdd AND2X2
XFILL_32_2_0 gnd vdd FILL
XDFFPOSX1_27 BUFX2_29/A CLKBUF1_1/Y AOI22X1_56/Y gnd vdd DFFPOSX1
XAOI21X1_328 INVX1_17/A AOI21X1_55/B BUFX4_92/Y gnd OAI21X1_794/C vdd AOI21X1
XAOI21X1_317 XNOR2X1_20/Y INVX1_298/Y BUFX4_27/Y gnd OAI21X1_757/C vdd AOI21X1
XAOI21X1_306 XNOR2X1_16/Y AOI21X1_51/B BUFX4_92/Y gnd OAI21X1_729/C vdd AOI21X1
XDFFPOSX1_16 BUFX2_18/A CLKBUF1_2/Y DFFPOSX1_16/D gnd vdd DFFPOSX1
XAOI21X1_339 XNOR2X1_6/Y OAI21X1_825/B BUFX4_96/Y gnd OAI21X1_825/C vdd AOI21X1
XDFFPOSX1_49 BUFX2_51/A CLKBUF1_4/Y DFFPOSX1_49/D gnd vdd DFFPOSX1
XDFFPOSX1_38 BUFX2_40/A CLKBUF1_8/Y AOI21X1_96/Y gnd vdd DFFPOSX1
XFILL_23_2_0 gnd vdd FILL
XFILL_6_3_0 gnd vdd FILL
XFILL_14_2_0 gnd vdd FILL
XINVX1_143 INVX1_143/A gnd INVX1_143/Y vdd INVX1
XINVX1_154 INVX1_154/A gnd INVX1_154/Y vdd INVX1
XINVX1_198 INVX1_198/A gnd INVX1_198/Y vdd INVX1
XINVX1_165 INVX1_165/A gnd INVX1_165/Y vdd INVX1
XINVX1_121 INVX1_121/A gnd INVX1_121/Y vdd INVX1
XINVX1_176 INVX1_176/A gnd INVX1_176/Y vdd INVX1
XINVX1_110 INVX1_110/A gnd INVX1_110/Y vdd INVX1
XINVX1_132 INVX1_132/A gnd INVX1_132/Y vdd INVX1
XINVX1_187 INVX1_187/A gnd INVX1_187/Y vdd INVX1
XNOR2X1_501 NOR2X1_501/A NOR2X1_501/B gnd NOR2X1_501/Y vdd NOR2X1
XAOI21X1_103 OR2X2_12/B OR2X2_12/A NOR2X1_173/Y gnd XNOR2X1_33/A vdd AOI21X1
XAOI21X1_114 INVX1_154/A INVX1_163/A BUFX4_93/Y gnd OAI21X1_363/C vdd AOI21X1
XAOI21X1_158 OAI21X1_453/Y AOI21X1_158/B NOR2X1_236/Y gnd DFFPOSX1_47/D vdd AOI21X1
XAOI21X1_125 INVX1_156/A INVX1_162/A NOR2X1_190/B gnd OAI21X1_424/A vdd AOI21X1
XAOI21X1_136 AOI21X1_136/A OR2X2_21/Y NAND3X1_20/Y gnd AOI21X1_137/B vdd AOI21X1
XAOI21X1_147 INVX4_21/A NOR2X1_226/Y BUFX4_27/Y gnd OAI21X1_437/C vdd AOI21X1
XAOI21X1_169 BUFX4_80/Y OAI21X1_483/Y OAI21X1_487/Y gnd AND2X2_28/A vdd AOI21X1
XFILL_30_5_1 gnd vdd FILL
XNAND2X1_309 BUFX4_134/Y INVX1_89/A gnd OAI21X1_291/C vdd NAND2X1
XNOR2X1_331 INVX2_84/Y AND2X2_41/A gnd NOR2X1_332/A vdd NOR2X1
XNOR2X1_320 NOR2X1_320/A NOR2X1_320/B gnd INVX2_82/A vdd NOR2X1
XNOR2X1_342 operand_A[60] operand_B[60] gnd NOR2X1_350/A vdd NOR2X1
XNOR2X1_386 BUFX2_53/A BUFX2_54/A gnd NOR2X1_386/Y vdd NOR2X1
XNOR2X1_353 BUFX4_98/Y BUFX2_63/A gnd NOR2X1_353/Y vdd NOR2X1
XNOR2X1_375 BUFX4_98/Y BUFX2_66/A gnd NOR2X1_375/Y vdd NOR2X1
XNOR2X1_364 operand_A[62] operand_B[62] gnd OAI22X1_22/D vdd NOR2X1
XFILL_21_5_1 gnd vdd FILL
XFILL_20_0_0 gnd vdd FILL
XOAI21X1_837 operand_A[12] operand_B[12] BUFX4_2/Y gnd OAI21X1_838/C vdd OAI21X1
XOAI21X1_804 AOI21X1_9/Y INVX1_17/A INVX1_305/Y gnd OAI21X1_805/B vdd OAI21X1
XNOR2X1_397 NOR2X1_397/A NOR2X1_397/B gnd NOR2X1_397/Y vdd NOR2X1
XOAI21X1_848 MUX2X1_64/S INVX1_328/A OAI21X1_848/C gnd AND2X2_62/A vdd OAI21X1
XOAI21X1_815 OAI21X1_815/A MUX2X1_34/S BUFX4_78/Y gnd OAI21X1_816/A vdd OAI21X1
XOAI21X1_826 INVX1_117/A BUFX4_24/Y OAI21X1_826/C gnd NOR2X1_461/B vdd OAI21X1
XOAI21X1_859 OAI21X1_859/A XNOR2X1_22/Y BUFX4_138/Y gnd OAI21X1_859/Y vdd OAI21X1
XFILL_28_1_0 gnd vdd FILL
XFILL_3_1_0 gnd vdd FILL
XFILL_12_5_1 gnd vdd FILL
XFILL_11_0_0 gnd vdd FILL
XFILL_19_1_0 gnd vdd FILL
XNOR2X1_82 NOR2X1_82/A NOR2X1_82/B gnd INVX1_52/A vdd NOR2X1
XNOR2X1_71 alu_op[1] INVX1_35/Y gnd INVX2_34/A vdd NOR2X1
XNAND3X1_71 NAND3X1_71/A NAND3X1_71/B OAI22X1_33/Y gnd NAND3X1_71/Y vdd NAND3X1
XNOR2X1_60 NOR2X1_60/A NOR2X1_60/B gnd NOR2X1_60/Y vdd NOR2X1
XNAND3X1_60 BUFX4_114/Y operand_A[5] BUFX4_150/Y gnd NAND3X1_61/B vdd NAND3X1
XNOR2X1_93 NOR2X1_93/A BUFX2_34/A gnd NOR2X1_93/Y vdd NOR2X1
XBUFX2_9 BUFX2_9/A gnd result[6] vdd BUFX2
XNAND2X1_139 INVX1_75/A AND2X2_6/A gnd OAI21X1_94/C vdd NAND2X1
XNAND2X1_4 operand_B[22] INVX4_3/Y gnd INVX1_3/A vdd NAND2X1
XNAND2X1_128 MUX2X1_87/S OAI21X1_76/Y gnd OAI21X1_79/C vdd NAND2X1
XNAND2X1_117 BUFX4_38/Y OR2X2_13/A gnd OAI21X1_74/C vdd NAND2X1
XNAND2X1_106 MUX2X1_9/S operand_A[7] gnd OAI21X1_57/C vdd NAND2X1
XNOR2X1_172 BUFX4_101/Y BUFX2_42/A gnd NOR2X1_172/Y vdd NOR2X1
XNOR2X1_183 NOR2X1_183/A NOR2X1_183/B gnd NOR2X1_184/B vdd NOR2X1
XNOR2X1_161 INVX1_72/Y BUFX4_8/Y gnd INVX1_145/A vdd NOR2X1
XNOR2X1_150 OR2X2_13/B MUX2X1_39/B gnd NOR2X1_150/Y vdd NOR2X1
XNOR2X1_194 MUX2X1_32/S OAI22X1_15/B gnd NOR2X1_194/Y vdd NOR2X1
XOAI21X1_601 INVX1_249/Y INVX1_240/Y OAI21X1_601/C gnd INVX1_253/A vdd OAI21X1
XOAI21X1_634 OAI22X1_9/C NOR2X1_371/A BUFX4_98/Y gnd NOR2X1_374/B vdd OAI21X1
XOAI21X1_667 NOR2X1_421/Y NOR2X1_183/B OAI21X1_667/C gnd OAI21X1_667/Y vdd OAI21X1
XOAI21X1_623 OAI21X1_623/A OR2X2_38/A INVX1_260/Y gnd OAI21X1_623/Y vdd OAI21X1
XOAI21X1_612 INVX1_257/A INVX1_255/A NOR2X1_359/A gnd OAI21X1_622/C vdd OAI21X1
XOAI21X1_656 INVX4_12/Y operand_B[61] OAI22X1_24/Y gnd OAI21X1_656/Y vdd OAI21X1
XOAI21X1_645 AND2X2_47/Y OAI21X1_645/B AND2X2_10/Y gnd AND2X2_48/A vdd OAI21X1
XINVX2_9 operand_A[1] gnd INVX2_9/Y vdd INVX2
XOAI21X1_689 INVX2_13/Y MUX2X1_9/S OAI21X1_57/C gnd MUX2X1_76/B vdd OAI21X1
XAOI21X1_9 OAI21X1_9/Y NOR2X1_24/Y AOI21X1_9/C gnd AOI21X1_9/Y vdd AOI21X1
XOAI21X1_678 MUX2X1_97/S MUX2X1_72/Y OAI21X1_678/C gnd MUX2X1_74/A vdd OAI21X1
XXNOR2X1_39 XNOR2X1_39/A INVX1_219/A gnd XNOR2X1_39/Y vdd XNOR2X1
XXNOR2X1_28 operand_A[25] operand_B[25] gnd XNOR2X1_47/B vdd XNOR2X1
XMUX2X1_112 MUX2X1_112/A OAI21X1_85/B BUFX4_16/Y gnd NOR2X1_446/B vdd MUX2X1
XXNOR2X1_17 BUFX4_35/Y operand_A[3] gnd XNOR2X1_17/Y vdd XNOR2X1
XMUX2X1_101 MUX2X1_114/B MUX2X1_113/A BUFX4_131/Y gnd MUX2X1_102/A vdd MUX2X1
XMUX2X1_123 MUX2X1_123/A MUX2X1_75/Y OR2X2_43/B gnd MUX2X1_123/Y vdd MUX2X1
XBUFX2_38 BUFX2_38/A gnd result[35] vdd BUFX2
XBUFX2_49 BUFX2_49/A gnd result[46] vdd BUFX2
XNAND2X1_651 NOR2X1_3/B OAI21X1_34/Y gnd OAI21X1_944/C vdd NAND2X1
XINVX1_63 INVX1_63/A gnd INVX1_63/Y vdd INVX1
XINVX1_41 INVX1_41/A gnd INVX1_41/Y vdd INVX1
XBUFX2_27 BUFX2_27/A gnd result[24] vdd BUFX2
XINVX1_74 INVX1_74/A gnd INVX1_74/Y vdd INVX1
XNAND2X1_640 AOI22X1_52/Y OAI22X1_32/Y gnd NAND2X1_640/Y vdd NAND2X1
XINVX1_52 INVX1_52/A gnd INVX1_52/Y vdd INVX1
XINVX1_96 INVX1_96/A gnd INVX1_96/Y vdd INVX1
XINVX1_85 INVX1_85/A gnd INVX1_85/Y vdd INVX1
XINVX1_30 INVX1_30/A gnd INVX1_30/Y vdd INVX1
XBUFX2_16 BUFX2_16/A gnd result[13] vdd BUFX2
XDFFPOSX1_4 BUFX2_6/A CLKBUF1_7/Y DFFPOSX1_4/D gnd vdd DFFPOSX1
XNOR2X1_7 INVX1_5/Y INVX4_6/Y gnd NOR2X1_7/Y vdd NOR2X1
XAOI21X1_39 AND2X2_6/Y NOR2X1_97/Y BUFX4_95/Y gnd AOI21X1_43/B vdd AOI21X1
XAOI21X1_17 NOR2X1_3/Y AND2X2_74/A INVX1_2/Y gnd INVX1_26/A vdd AOI21X1
XAOI21X1_28 NOR2X1_30/Y XNOR2X1_6/Y INVX1_83/A gnd OAI21X1_30/C vdd AOI21X1
XFILL_26_4_1 gnd vdd FILL
XOAI22X1_25 INVX1_230/Y operand_A[56] operand_A[57] INVX1_235/Y gnd OAI22X1_25/Y vdd
+ OAI22X1
XOAI22X1_36 OAI22X1_36/A OAI22X1_36/B OAI22X1_36/C OAI22X1_36/D gnd OAI22X1_36/Y vdd
+ OAI22X1
XOAI22X1_14 INVX2_49/Y INVX1_151/A OAI22X1_14/C BUFX4_10/Y gnd OAI22X1_33/B vdd OAI22X1
XFILL_1_4_1 gnd vdd FILL
XOAI21X1_486 BUFX4_61/Y INVX1_201/Y AOI22X1_18/Y gnd NOR2X1_254/B vdd OAI21X1
XOAI21X1_453 INVX1_186/A OAI21X1_453/B OAI21X1_453/C gnd OAI21X1_453/Y vdd OAI21X1
XOAI21X1_475 NOR2X1_231/B NOR2X1_231/A INVX4_22/A gnd OR2X2_29/B vdd OAI21X1
XOAI21X1_464 operand_A[47] operand_B[47] BUFX4_5/Y gnd NAND3X1_28/A vdd OAI21X1
XOAI21X1_442 INVX1_165/Y BUFX4_120/Y OAI21X1_442/C gnd INVX1_181/A vdd OAI21X1
XOAI21X1_497 BUFX4_111/Y AOI22X1_19/Y OAI21X1_497/C gnd OAI21X1_497/Y vdd OAI21X1
XOAI21X1_420 NOR2X1_80/A OAI22X1_18/B OAI21X1_420/C gnd AND2X2_59/A vdd OAI21X1
XOAI21X1_431 BUFX4_23/Y MUX2X1_31/A OAI21X1_431/C gnd OAI21X1_435/B vdd OAI21X1
XNAND2X1_470 BUFX4_43/Y operand_A[52] gnd OAI21X1_534/C vdd NAND2X1
XNAND2X1_481 BUFX4_70/Y OAI21X1_577/B gnd OAI21X1_557/C vdd NAND2X1
XFILL_8_0_0 gnd vdd FILL
XFILL_9_5_1 gnd vdd FILL
XNAND2X1_492 NAND2X1_492/A NAND2X1_492/B gnd NOR2X1_314/A vdd NAND2X1
XFILL_17_4_1 gnd vdd FILL
XOAI21X1_80 INVX2_46/Y MUX2X1_4/S OAI21X1_80/C gnd OAI21X1_80/Y vdd OAI21X1
XOAI21X1_91 INVX1_56/Y INVX2_49/Y BUFX4_114/Y gnd OAI22X1_2/B vdd OAI21X1
XOAI21X1_250 AOI21X1_71/Y BUFX4_16/Y OAI21X1_251/C gnd OAI21X1_250/Y vdd OAI21X1
XOAI21X1_283 INVX2_62/A INVX4_17/A OAI21X1_283/C gnd AOI21X1_82/C vdd OAI21X1
XAND2X2_50 AND2X2_50/A AND2X2_50/B gnd AND2X2_50/Y vdd AND2X2
XINVX1_325 INVX1_325/A gnd INVX1_325/Y vdd INVX1
XOAI21X1_294 INVX1_130/Y MUX2X1_98/S OAI21X1_294/C gnd INVX1_131/A vdd OAI21X1
XOAI21X1_272 OAI21X1_272/A XOR2X1_7/A INVX1_118/Y gnd AND2X2_20/A vdd OAI21X1
XAND2X2_72 AND2X2_72/A OR2X2_48/Y gnd AND2X2_72/Y vdd AND2X2
XINVX1_314 INVX1_314/A gnd INVX1_314/Y vdd INVX1
XINVX1_303 NOR2X1_26/Y gnd INVX1_303/Y vdd INVX1
XOAI21X1_261 MUX2X1_32/S OAI21X1_261/B OAI21X1_261/C gnd AOI21X1_74/B vdd OAI21X1
XAND2X2_61 AND2X2_61/A AND2X2_61/B gnd AND2X2_61/Y vdd AND2X2
XFILL_32_2_1 gnd vdd FILL
XAOI21X1_307 XNOR2X1_16/Y OAI21X1_9/A BUFX4_27/Y gnd AOI21X1_308/B vdd AOI21X1
XDFFPOSX1_39 OR2X2_36/A CLKBUF1_3/Y OAI21X1_345/Y gnd vdd DFFPOSX1
XDFFPOSX1_28 BUFX2_30/A CLKBUF1_1/Y AOI22X1_57/Y gnd vdd DFFPOSX1
XAOI21X1_318 XNOR2X1_20/Y OAI21X1_759/B BUFX4_92/Y gnd OAI21X1_759/C vdd AOI21X1
XAOI21X1_329 OR2X2_13/B MUX2X1_75/A BUFX4_186/Y gnd OAI21X1_796/C vdd AOI21X1
XDFFPOSX1_17 BUFX2_19/A CLKBUF1_2/Y AOI22X1_45/Y gnd vdd DFFPOSX1
XFILL_23_2_1 gnd vdd FILL
XFILL_6_3_1 gnd vdd FILL
XFILL_14_2_1 gnd vdd FILL
XINVX1_100 INVX1_100/A gnd INVX1_100/Y vdd INVX1
XINVX1_144 INVX1_144/A gnd INVX1_144/Y vdd INVX1
XINVX1_155 INVX1_155/A gnd INVX1_155/Y vdd INVX1
XINVX1_199 INVX1_199/A gnd INVX1_199/Y vdd INVX1
XINVX1_188 INVX1_188/A gnd INVX1_188/Y vdd INVX1
XINVX1_133 INVX1_133/A gnd INVX1_133/Y vdd INVX1
XINVX1_111 INVX1_111/A gnd INVX1_111/Y vdd INVX1
XINVX1_122 INVX1_122/A gnd INVX1_122/Y vdd INVX1
XINVX1_166 NAND3X1_7/C gnd INVX1_166/Y vdd INVX1
XINVX1_177 INVX1_177/A gnd INVX1_177/Y vdd INVX1
XNOR2X1_502 BUFX4_9/Y OAI22X1_18/C gnd OAI22X1_37/A vdd NOR2X1
XAOI21X1_104 BUFX4_5/Y NAND2X1_355/B NOR2X1_174/Y gnd OAI21X1_354/C vdd AOI21X1
XAOI21X1_126 INVX1_169/A OAI21X1_393/B BUFX4_30/Y gnd OAI21X1_393/C vdd AOI21X1
XFILL_27_1 gnd vdd FILL
XAOI21X1_137 OAI21X1_409/Y AOI21X1_137/B NOR2X1_214/Y gnd DFFPOSX1_44/D vdd AOI21X1
XAOI21X1_115 NAND2X1_362/Y AOI21X1_115/B OAI21X1_364/Y gnd AND2X2_15/A vdd AOI21X1
XAOI21X1_148 BUFX4_163/Y NOR2X1_361/B INVX8_15/Y gnd NAND2X1_417/B vdd AOI21X1
XAOI21X1_159 INVX1_186/A OAI21X1_453/B NOR2X1_231/B gnd XNOR2X1_35/A vdd AOI21X1
XNOR2X1_376 BUFX2_39/A BUFX2_40/A gnd NOR2X1_376/Y vdd NOR2X1
XNOR2X1_310 INVX2_79/A INVX1_224/A gnd NOR2X1_310/Y vdd NOR2X1
XNOR2X1_332 NOR2X1_332/A AND2X2_41/Y gnd NOR2X1_332/Y vdd NOR2X1
XNOR2X1_321 NOR2X1_321/A NOR2X1_321/B gnd NOR2X1_321/Y vdd NOR2X1
XNOR2X1_365 INVX2_90/Y INVX1_256/Y gnd INVX2_91/A vdd NOR2X1
XNOR2X1_343 INVX2_87/Y INVX1_245/Y gnd INVX1_251/A vdd NOR2X1
XNOR2X1_354 INVX4_12/Y INVX1_252/Y gnd INVX1_257/A vdd NOR2X1
XNOR2X1_387 BUFX2_51/A BUFX2_52/A gnd NOR2X1_387/Y vdd NOR2X1
XFILL_20_0_1 gnd vdd FILL
XOAI21X1_838 BUFX4_154/Y XNOR2X1_5/Y OAI21X1_838/C gnd NOR2X1_468/A vdd OAI21X1
XOAI21X1_805 INVX2_17/Y OAI21X1_805/B OAI21X1_805/C gnd AOI22X1_39/D vdd OAI21X1
XOAI21X1_827 BUFX4_37/Y MUX2X1_102/A OAI21X1_827/C gnd OAI21X1_828/A vdd OAI21X1
XNOR2X1_398 BUFX2_6/A BUFX2_5/A gnd NOR2X1_398/Y vdd NOR2X1
XOAI21X1_816 OAI21X1_816/A NOR2X1_458/Y INVX8_9/A gnd OAI21X1_817/C vdd OAI21X1
XOAI21X1_849 AND2X2_62/Y AND2X2_63/Y BUFX4_89/Y gnd NAND3X1_66/B vdd OAI21X1
XFILL_28_1_1 gnd vdd FILL
XFILL_3_1_1 gnd vdd FILL
XFILL_11_0_1 gnd vdd FILL
XNAND3X1_50 INVX1_274/Y INVX1_275/Y NOR2X1_404/Y gnd NOR2X1_406/A vdd NAND3X1
XNOR2X1_94 AND2X2_5/Y NOR2X1_94/B gnd NOR2X1_94/Y vdd NOR2X1
XNAND3X1_72 NAND3X1_72/A NAND3X1_72/B OAI22X1_34/Y gnd NOR2X1_499/B vdd NAND3X1
XFILL_19_1_1 gnd vdd FILL
XNOR2X1_72 INVX2_33/Y INVX2_34/Y gnd NOR2X1_72/Y vdd NOR2X1
XNOR2X1_83 NOR2X1_83/A INVX1_52/Y gnd INVX1_55/A vdd NOR2X1
XNOR2X1_61 operand_B[9] INVX2_24/Y gnd NOR2X1_61/Y vdd NOR2X1
XNAND3X1_61 NAND3X1_61/A NAND3X1_61/B NAND3X1_61/C gnd NAND3X1_61/Y vdd NAND3X1
XNOR2X1_50 operand_B[18] INVX4_5/Y gnd NOR2X1_50/Y vdd NOR2X1
XNAND2X1_107 MUX2X1_97/S OAI21X1_57/Y gnd OAI21X1_58/C vdd NAND2X1
XNAND2X1_129 BUFX4_53/Y operand_A[33] gnd OAI21X1_77/C vdd NAND2X1
XNAND2X1_118 MUX2X1_3/S operand_A[53] gnd OAI21X1_67/C vdd NAND2X1
XNAND2X1_5 operand_B[21] INVX4_4/Y gnd INVX1_4/A vdd NAND2X1
XNOR2X1_173 operand_B[38] INVX2_66/Y gnd NOR2X1_173/Y vdd NOR2X1
XNOR2X1_184 NOR2X1_184/A NOR2X1_184/B gnd AND2X2_27/A vdd NOR2X1
XNOR2X1_162 OAI22X1_4/Y NOR2X1_162/B gnd NOR2X1_162/Y vdd NOR2X1
XNOR2X1_140 BUFX4_113/Y BUFX4_171/Y gnd INVX8_18/A vdd NOR2X1
XNOR2X1_151 INVX4_10/Y MUX2X1_71/S gnd INVX1_118/A vdd NOR2X1
XMUX2X1_90 MUX2X1_90/A MUX2X1_90/B BUFX4_66/Y gnd MUX2X1_94/B vdd MUX2X1
XNOR2X1_195 MUX2X1_34/S OAI22X1_15/C gnd NOR2X1_195/Y vdd NOR2X1
XOAI21X1_657 INVX4_13/Y operand_B[57] OAI22X1_25/Y gnd OAI21X1_658/B vdd OAI21X1
XOAI21X1_635 BUFX4_157/Y INVX4_25/Y OAI21X1_635/C gnd NOR2X1_374/A vdd OAI21X1
XOAI21X1_602 OAI21X1_623/A INVX2_88/A BUFX4_143/Y gnd OAI21X1_602/Y vdd OAI21X1
XOAI21X1_624 INVX2_90/Y BUFX4_43/Y OAI21X1_624/C gnd MUX2X1_65/A vdd OAI21X1
XOAI21X1_668 NOR2X1_250/Y NOR2X1_422/Y OAI21X1_668/C gnd OAI21X1_673/C vdd OAI21X1
XOAI21X1_613 INVX4_12/Y MUX2X1_3/S OAI21X1_613/C gnd INVX1_254/A vdd OAI21X1
XOAI21X1_646 NOR2X1_53/Y INVX1_3/A NAND2X1_65/Y gnd OAI21X1_651/B vdd OAI21X1
XOAI21X1_679 INVX2_6/Y BUFX4_50/Y OAI21X1_37/C gnd INVX1_285/A vdd OAI21X1
XMUX2X1_113 MUX2X1_113/A MUX2X1_99/A INVX8_3/A gnd MUX2X1_115/B vdd MUX2X1
XMUX2X1_102 MUX2X1_102/A MUX2X1_99/Y XOR2X1_4/A gnd MUX2X1_102/Y vdd MUX2X1
XNAND2X1_641 OAI21X1_902/Y NAND2X1_641/B gnd OAI21X1_904/A vdd NAND2X1
XXNOR2X1_29 operand_A[24] operand_B[24] gnd XNOR2X1_29/Y vdd XNOR2X1
XINVX1_31 INVX1_31/A gnd INVX1_31/Y vdd INVX1
XINVX1_20 operand_B[8] gnd INVX1_20/Y vdd INVX1
XXNOR2X1_18 operand_B[7] operand_A[7] gnd XNOR2X1_18/Y vdd XNOR2X1
XMUX2X1_124 MUX2X1_124/A MUX2X1_124/B BUFX4_162/Y gnd MUX2X1_124/Y vdd MUX2X1
XINVX1_42 INVX1_42/A gnd INVX1_42/Y vdd INVX1
XNAND2X1_630 OR2X2_7/B NOR2X1_145/B gnd OAI21X1_882/C vdd NAND2X1
XBUFX2_39 BUFX2_39/A gnd result[36] vdd BUFX2
XINVX1_75 INVX1_75/A gnd INVX1_75/Y vdd INVX1
XINVX1_97 INVX1_97/A gnd INVX1_97/Y vdd INVX1
XBUFX2_28 BUFX2_28/A gnd result[25] vdd BUFX2
XINVX1_53 INVX1_53/A gnd INVX1_53/Y vdd INVX1
XDFFPOSX1_5 BUFX2_7/A CLKBUF1_7/Y DFFPOSX1_5/D gnd vdd DFFPOSX1
XBUFX2_17 BUFX2_17/A gnd result[14] vdd BUFX2
XINVX1_64 INVX1_64/A gnd INVX1_64/Y vdd INVX1
XINVX1_86 INVX1_86/A gnd INVX1_86/Y vdd INVX1
XNOR2X1_8 INVX1_6/Y INVX2_6/Y gnd OR2X2_46/B vdd NOR2X1
XAOI21X1_29 NAND2X1_36/B NOR2X1_65/Y NOR2X1_64/Y gnd INVX1_84/A vdd AOI21X1
XAOI21X1_18 INVX1_11/A NOR2X1_49/Y OAI21X1_7/B gnd INVX1_316/A vdd AOI21X1
XOAI22X1_26 INVX2_76/Y operand_A[50] operand_A[51] INVX2_77/Y gnd OAI22X1_26/Y vdd
+ OAI22X1
XOAI21X1_410 INVX2_71/Y operand_B[42] AND2X2_19/A gnd OR2X2_21/A vdd OAI21X1
XOAI21X1_421 INVX2_73/Y operand_B[43] NAND3X1_21/Y gnd OAI21X1_421/Y vdd OAI21X1
XOAI21X1_432 INVX2_46/Y MUX2X1_9/S OAI21X1_432/C gnd OAI21X1_457/B vdd OAI21X1
XOAI22X1_37 OAI22X1_37/A OAI22X1_37/B OAI22X1_37/C OAI22X1_37/D gnd OAI22X1_37/Y vdd
+ OAI22X1
XOAI22X1_15 INVX8_8/Y OAI22X1_15/B OAI22X1_15/C OAI22X1_1/B gnd OAI22X1_35/D vdd OAI22X1
XOAI21X1_498 INVX4_23/Y NOR2X1_272/B OAI21X1_498/C gnd OAI21X1_498/Y vdd OAI21X1
XOAI21X1_476 INVX1_192/Y NOR2X1_250/Y OAI21X1_668/C gnd OR2X2_30/B vdd OAI21X1
XOAI21X1_454 OAI21X1_454/A INVX4_21/Y NOR2X1_249/B gnd OR2X2_24/A vdd OAI21X1
XOAI21X1_487 NOR2X1_484/B OR2X2_32/B NOR2X1_254/Y gnd OAI21X1_487/Y vdd OAI21X1
XOAI21X1_465 OR2X2_25/B NOR2X1_478/B OAI21X1_465/C gnd OR2X2_27/A vdd OAI21X1
XOAI21X1_443 BUFX4_25/Y OAI21X1_443/B OAI21X1_443/C gnd NOR2X1_361/B vdd OAI21X1
XNAND2X1_460 INVX4_23/A INVX1_212/A gnd NOR2X1_278/B vdd NAND2X1
XNAND2X1_471 NOR2X1_82/A OAI21X1_511/Y gnd OAI21X1_535/C vdd NAND2X1
XNAND2X1_493 BUFX4_133/Y OAI21X1_526/Y gnd OAI21X1_568/C vdd NAND2X1
XNAND2X1_482 MUX2X1_62/S INVX1_227/Y gnd OAI21X1_558/C vdd NAND2X1
XFILL_8_0_1 gnd vdd FILL
XOAI21X1_70 INVX2_42/Y BUFX4_46/Y OAI21X1_70/C gnd INVX1_49/A vdd OAI21X1
XOAI21X1_81 BUFX4_192/Y MUX2X1_8/Y OAI21X1_81/C gnd INVX1_50/A vdd OAI21X1
XOAI21X1_92 operand_A[30] operand_B[30] BUFX4_6/Y gnd AND2X2_4/A vdd OAI21X1
XOAI21X1_240 INVX1_77/A OAI21X1_240/B INVX1_108/Y gnd AND2X2_12/A vdd OAI21X1
XOAI21X1_251 BUFX4_16/Y INVX1_109/Y OAI21X1_251/C gnd INVX1_110/A vdd OAI21X1
XOAI21X1_262 OR2X2_25/B INVX1_111/Y AOI21X1_74/Y gnd AOI21X1_75/C vdd OAI21X1
XOAI21X1_273 BUFX4_179/Y NOR2X1_145/B OAI21X1_273/C gnd AOI22X1_7/C vdd OAI21X1
XOAI21X1_284 INVX1_77/A OR2X2_17/A AOI21X1_82/Y gnd INVX2_64/A vdd OAI21X1
XINVX1_326 NOR2X1_3/B gnd INVX1_326/Y vdd INVX1
XAND2X2_40 INVX8_13/Y AND2X2_40/B gnd AND2X2_40/Y vdd AND2X2
XAND2X2_73 AND2X2_73/A INVX2_94/Y gnd OR2X2_49/A vdd AND2X2
XOAI21X1_295 INVX1_131/Y XOR2X1_7/A OAI21X1_295/C gnd MUX2X1_40/B vdd OAI21X1
XAND2X2_51 AND2X2_51/A AND2X2_51/B gnd AND2X2_51/Y vdd AND2X2
XINVX1_304 BUFX2_10/A gnd INVX1_304/Y vdd INVX1
XAND2X2_62 AND2X2_62/A BUFX4_82/Y gnd AND2X2_62/Y vdd AND2X2
XINVX1_315 INVX1_315/A gnd INVX1_315/Y vdd INVX1
XNAND2X1_290 MUX2X1_99/S INVX1_69/Y gnd OAI21X1_265/C vdd NAND2X1
XAOI21X1_308 OAI21X1_741/C AOI21X1_308/B NAND3X1_57/Y gnd NAND3X1_58/B vdd AOI21X1
XAOI21X1_319 BUFX4_162/Y MUX2X1_109/Y NOR2X1_442/Y gnd OR2X2_40/A vdd AOI21X1
XDFFPOSX1_29 BUFX2_31/A CLKBUF1_1/Y DFFPOSX1_29/D gnd vdd DFFPOSX1
XDFFPOSX1_18 BUFX2_20/A CLKBUF1_2/Y AOI22X1_47/Y gnd vdd DFFPOSX1
XINVX1_134 INVX1_134/A gnd INVX1_134/Y vdd INVX1
XINVX1_101 INVX1_101/A gnd INVX1_101/Y vdd INVX1
XINVX1_123 INVX1_123/A gnd INVX1_123/Y vdd INVX1
XINVX1_112 INVX1_112/A gnd INVX1_112/Y vdd INVX1
XINVX1_156 INVX1_156/A gnd INVX1_156/Y vdd INVX1
XINVX1_178 INVX1_178/A gnd INVX1_178/Y vdd INVX1
XINVX1_145 INVX1_145/A gnd INVX1_145/Y vdd INVX1
XINVX1_189 INVX1_189/A gnd INVX1_189/Y vdd INVX1
XINVX1_167 MUX2X1_29/B gnd INVX1_167/Y vdd INVX1
XNOR2X1_503 NOR2X1_503/A NOR2X1_503/B gnd NOR2X1_503/Y vdd NOR2X1
XFILL_27_2 gnd vdd FILL
XAOI21X1_138 NOR2X1_218/Y NOR2X1_203/A OAI21X1_421/Y gnd NOR2X1_248/B vdd AOI21X1
XAOI21X1_127 MUX2X1_57/S OAI21X1_406/Y NOR2X1_205/Y gnd OR2X2_19/A vdd AOI21X1
XAOI21X1_116 BUFX4_186/Y INVX2_48/A AND2X2_57/A gnd NOR2X1_452/B vdd AOI21X1
XAOI21X1_105 BUFX4_84/Y OAI21X1_353/Y OAI21X1_355/Y gnd NAND3X1_15/B vdd AOI21X1
XAOI21X1_149 INVX4_18/A NOR2X1_227/Y NAND3X1_23/Y gnd NAND3X1_24/A vdd AOI21X1
XFILL_24_5_0 gnd vdd FILL
XINVX4_20 INVX4_20/A gnd OR2X2_19/B vdd INVX4
XFILL_15_5_0 gnd vdd FILL
XNOR2X1_388 BUFX2_49/A BUFX2_50/A gnd NOR2X1_388/Y vdd NOR2X1
XNOR2X1_377 BUFX2_37/A BUFX2_38/A gnd NOR2X1_377/Y vdd NOR2X1
XNOR2X1_311 NOR2X1_312/A NOR2X1_311/B gnd INVX1_233/A vdd NOR2X1
XNOR2X1_399 BUFX2_65/A BUFX2_66/A gnd NOR2X1_399/Y vdd NOR2X1
XNOR2X1_333 NOR2X1_333/A BUFX4_145/Y gnd NOR2X1_334/A vdd NOR2X1
XNOR2X1_366 INVX2_88/Y INVX4_24/Y gnd INVX1_258/A vdd NOR2X1
XNOR2X1_322 operand_B[56] INVX2_39/Y gnd NOR2X1_323/A vdd NOR2X1
XNOR2X1_344 NOR2X1_350/A INVX1_251/A gnd INVX2_88/A vdd NOR2X1
XNOR2X1_355 operand_A[61] operand_B[61] gnd INVX1_255/A vdd NOR2X1
XNOR2X1_300 MUX2X1_25/S NOR2X1_300/B gnd NOR2X1_301/A vdd NOR2X1
XOAI21X1_806 OAI21X1_32/A INVX1_278/Y OAI21X1_806/C gnd OAI21X1_807/A vdd OAI21X1
XOAI21X1_828 OAI21X1_828/A OR2X2_7/B BUFX4_78/Y gnd NOR2X1_462/B vdd OAI21X1
XOAI21X1_817 INVX8_8/Y OAI22X1_16/A OAI21X1_817/C gnd OAI21X1_817/Y vdd OAI21X1
XOAI21X1_839 NOR2X1_467/Y NOR2X1_466/Y INVX8_10/A gnd OAI21X1_840/C vdd OAI21X1
XNAND3X1_40 INVX4_25/A NAND3X1_40/B NAND3X1_40/C gnd NAND3X1_40/Y vdd NAND3X1
XNAND3X1_51 INVX1_276/Y INVX1_277/Y NOR2X1_405/Y gnd NOR2X1_406/B vdd NAND3X1
XNAND3X1_62 NAND3X1_62/A NAND3X1_62/B NAND3X1_62/C gnd NAND3X1_62/Y vdd NAND3X1
XNOR2X1_95 operand_B[30] INVX2_35/Y gnd NOR2X1_97/A vdd NOR2X1
XNOR2X1_73 alu_op[3] INVX1_43/Y gnd INVX2_36/A vdd NOR2X1
XNOR2X1_84 INVX8_2/A INVX1_55/Y gnd INVX1_56/A vdd NOR2X1
XNOR2X1_62 operand_B[8] INVX2_26/Y gnd NOR2X1_62/Y vdd NOR2X1
XNOR2X1_40 INVX1_16/Y INVX2_16/Y gnd NOR2X1_40/Y vdd NOR2X1
XNOR2X1_51 operand_B[19] INVX2_7/Y gnd NOR2X1_51/Y vdd NOR2X1
XFILL_30_3_0 gnd vdd FILL
XNAND2X1_119 BUFX4_43/Y operand_A[51] gnd OAI21X1_68/C vdd NAND2X1
XNAND2X1_108 BUFX4_131/Y OAI21X1_58/Y gnd OAI21X1_59/C vdd NAND2X1
XNAND2X1_6 operand_A[20] INVX2_3/Y gnd NAND2X1_8/A vdd NAND2X1
XNOR2X1_152 NOR2X1_93/A BUFX2_38/A gnd NOR2X1_152/Y vdd NOR2X1
XNOR2X1_163 BUFX4_101/Y BUFX2_40/A gnd NOR2X1_163/Y vdd NOR2X1
XNOR2X1_174 NOR2X1_174/A BUFX4_61/Y gnd NOR2X1_174/Y vdd NOR2X1
XNOR2X1_130 BUFX4_99/Y BUFX2_35/A gnd NOR2X1_130/Y vdd NOR2X1
XNOR2X1_185 NOR2X1_185/A OAI22X1_9/C gnd NOR2X1_185/Y vdd NOR2X1
XFILL_21_3_0 gnd vdd FILL
XOAI21X1_614 BUFX4_70/Y OAI21X1_614/B OAI21X1_614/C gnd MUX2X1_62/A vdd OAI21X1
XOAI21X1_603 INVX1_176/A INVX1_250/Y BUFX4_159/Y gnd OAI21X1_603/Y vdd OAI21X1
XNOR2X1_196 OR2X2_19/B NOR2X1_196/B gnd NOR2X1_199/A vdd NOR2X1
XMUX2X1_91 operand_A[12] operand_A[11] MUX2X1_1/S gnd MUX2X1_93/B vdd MUX2X1
XNOR2X1_141 NOR2X1_83/A MUX2X1_2/B gnd NOR2X1_141/Y vdd NOR2X1
XMUX2X1_80 operand_A[20] operand_A[19] MUX2X1_3/S gnd MUX2X1_80/Y vdd MUX2X1
XOAI21X1_658 INVX1_249/Y OAI21X1_658/B OAI21X1_658/C gnd OAI21X1_663/B vdd OAI21X1
XOAI21X1_669 INVX4_21/Y OAI21X1_669/B OAI21X1_669/C gnd NOR2X1_423/A vdd OAI21X1
XMUX2X1_103 MUX2X1_24/A MUX2X1_71/B MUX2X1_51/S gnd MUX2X1_121/B vdd MUX2X1
XOAI21X1_636 INVX1_51/A alu_op[2] alu_op[3] gnd DFFSR_1/D vdd OAI21X1
XOAI21X1_625 MUX2X1_67/Y INVX8_8/Y OAI21X1_625/C gnd OAI22X1_21/B vdd OAI21X1
XMUX2X1_125 AND2X2_14/A NOR2X1_446/B BUFX4_183/Y gnd MUX2X1_125/Y vdd MUX2X1
XMUX2X1_114 MUX2X1_114/A MUX2X1_114/B NOR2X1_83/A gnd MUX2X1_122/B vdd MUX2X1
XOAI21X1_647 OAI21X1_7/B NAND2X1_19/B INVX1_11/A gnd OAI21X1_647/Y vdd OAI21X1
XNAND2X1_642 INVX2_94/A OAI21X1_902/B gnd OAI21X1_906/C vdd NAND2X1
XINVX1_76 INVX1_76/A gnd INVX1_76/Y vdd INVX1
XINVX1_32 INVX1_32/A gnd INVX1_32/Y vdd INVX1
XINVX1_10 INVX1_10/A gnd INVX1_10/Y vdd INVX1
XINVX1_43 alu_op[2] gnd INVX1_43/Y vdd INVX1
XINVX1_54 INVX1_54/A gnd INVX1_54/Y vdd INVX1
XINVX1_65 INVX1_65/A gnd INVX1_65/Y vdd INVX1
XINVX1_21 INVX1_21/A gnd INVX1_21/Y vdd INVX1
XXNOR2X1_19 operand_A[6] operand_B[6] gnd XNOR2X1_19/Y vdd XNOR2X1
XNAND2X1_631 NOR2X1_490/Y OAI22X1_30/Y gnd NAND2X1_631/Y vdd NAND2X1
XNAND2X1_620 NOR2X1_75/A MUX2X1_129/B gnd AND2X2_61/B vdd NAND2X1
XFILL_29_4_0 gnd vdd FILL
XBUFX2_29 BUFX2_29/A gnd result[26] vdd BUFX2
XINVX1_87 INVX1_87/A gnd INVX1_87/Y vdd INVX1
XFILL_4_4_0 gnd vdd FILL
XINVX1_98 INVX1_98/A gnd INVX1_98/Y vdd INVX1
XDFFPOSX1_6 BUFX2_8/A CLKBUF1_7/Y DFFPOSX1_6/D gnd vdd DFFPOSX1
XBUFX2_18 BUFX2_18/A gnd result[15] vdd BUFX2
XFILL_12_3_0 gnd vdd FILL
XNOR2X1_9 INVX1_7/Y INVX2_7/Y gnd NOR2X1_9/Y vdd NOR2X1
XAOI21X1_19 NAND2X1_63/Y NOR2X1_50/Y NOR2X1_51/Y gnd OAI21X1_26/C vdd AOI21X1
XOAI21X1_422 INVX1_163/A NOR2X1_247/B NOR2X1_248/B gnd OAI21X1_423/B vdd OAI21X1
XOAI21X1_400 INVX2_71/Y MUX2X1_8/S OAI21X1_82/C gnd INVX1_171/A vdd OAI21X1
XOAI21X1_433 INVX1_171/Y BUFX4_73/Y OAI21X1_433/C gnd INVX1_178/A vdd OAI21X1
XOAI22X1_38 OAI22X1_38/A OAI22X1_38/B AND2X2_75/Y OAI22X1_38/D gnd OAI22X1_38/Y vdd
+ OAI22X1
XOAI22X1_27 OAI22X1_27/A OAI22X1_27/B OAI22X1_27/C AND2X2_55/Y gnd OAI22X1_27/Y vdd
+ OAI22X1
XOAI21X1_466 MUX2X1_21/A BUFX4_183/Y INVX4_11/Y gnd INVX1_195/A vdd OAI21X1
XOAI22X1_16 OAI22X1_16/A OAI22X1_1/B INVX1_170/Y INVX8_8/Y gnd OAI22X1_36/D vdd OAI22X1
XOAI21X1_444 MUX2X1_35/Y BUFX4_37/Y OAI21X1_444/C gnd MUX2X1_64/B vdd OAI21X1
XOAI21X1_411 BUFX4_20/Y OAI21X1_411/B OAI21X1_411/C gnd OAI22X1_19/C vdd OAI21X1
XOAI21X1_455 OAI22X1_1/A INVX8_8/Y INVX8_15/Y gnd OAI21X1_460/C vdd OAI21X1
XOAI21X1_488 INVX1_204/Y NOR2X1_259/Y OAI21X1_488/C gnd OAI21X1_488/Y vdd OAI21X1
XOAI21X1_477 AND2X2_27/Y INVX1_200/Y NOR2X1_251/Y gnd OAI21X1_477/Y vdd OAI21X1
XOAI21X1_499 NOR2X1_248/B OR2X2_29/Y NOR2X1_264/Y gnd OAI21X1_499/Y vdd OAI21X1
XNAND2X1_450 operand_A[49] INVX1_203/Y gnd OAI21X1_501/C vdd NAND2X1
XNAND2X1_461 operand_A[51] INVX2_77/Y gnd AOI22X1_30/A vdd NAND2X1
XNAND2X1_472 MUX2X1_66/S OAI21X1_535/Y gnd OAI21X1_536/C vdd NAND2X1
XNAND2X1_494 NAND2X1_494/A OAI21X1_569/Y gnd NAND2X1_494/Y vdd NAND2X1
XNAND2X1_483 BUFX4_36/Y OAI21X1_469/Y gnd OAI21X1_559/C vdd NAND2X1
XFILL_8_1 gnd vdd FILL
XOAI21X1_93 OAI21X1_94/C NOR2X1_94/Y OAI21X1_93/C gnd OAI21X1_93/Y vdd OAI21X1
XOAI21X1_82 INVX2_47/Y MUX2X1_5/S OAI21X1_82/C gnd OAI21X1_82/Y vdd OAI21X1
XOAI21X1_71 INVX2_43/Y BUFX4_48/Y OAI21X1_71/C gnd INVX1_87/A vdd OAI21X1
XOAI21X1_60 MUX2X1_2/Y BUFX4_20/Y OAI21X1_60/C gnd OAI22X1_1/A vdd OAI21X1
XFILL_26_2_0 gnd vdd FILL
XFILL_1_2_0 gnd vdd FILL
XOAI21X1_263 INVX2_62/A NOR2X1_144/Y AOI21X1_77/Y gnd AOI21X1_81/A vdd OAI21X1
XOAI21X1_241 INVX2_59/A AND2X2_12/A NOR2X1_136/Y gnd AOI21X1_76/A vdd OAI21X1
XOAI21X1_285 INVX2_64/Y INVX4_19/Y BUFX4_107/Y gnd AOI21X1_83/C vdd OAI21X1
XOAI21X1_230 BUFX4_68/Y MUX2X1_16/Y OAI21X1_230/C gnd OAI21X1_308/B vdd OAI21X1
XOAI21X1_252 INVX1_110/Y BUFX4_159/Y AOI21X1_72/A gnd INVX1_111/A vdd OAI21X1
XINVX1_305 NOR2X1_33/Y gnd INVX1_305/Y vdd INVX1
XOAI21X1_274 INVX1_62/Y NOR2X1_83/A OAI21X1_274/C gnd INVX1_120/A vdd OAI21X1
XOAI21X1_296 INVX1_129/Y BUFX4_19/Y OAI21X1_296/C gnd MUX2X1_32/A vdd OAI21X1
XINVX1_316 INVX1_316/A gnd INVX1_316/Y vdd INVX1
XAND2X2_41 AND2X2_41/A INVX2_84/Y gnd AND2X2_41/Y vdd AND2X2
XAND2X2_74 AND2X2_74/A INVX1_326/Y gnd AND2X2_74/Y vdd AND2X2
XINVX1_327 NOR2X1_2/Y gnd INVX1_327/Y vdd INVX1
XAND2X2_30 INVX8_13/Y AND2X2_30/B gnd AND2X2_30/Y vdd AND2X2
XAND2X2_52 AND2X2_52/A BUFX4_91/Y gnd AND2X2_52/Y vdd AND2X2
XFILL_9_3_0 gnd vdd FILL
XAND2X2_63 AND2X2_63/A BUFX4_111/Y gnd AND2X2_63/Y vdd AND2X2
XFILL_17_2_0 gnd vdd FILL
XNAND2X1_291 BUFX4_36/Y MUX2X1_39/A gnd OAI21X1_267/C vdd NAND2X1
XNAND2X1_280 BUFX4_119/Y INVX1_40/A gnd OAI21X1_256/C vdd NAND2X1
XAOI21X1_309 NOR2X1_433/Y OAI21X1_715/Y NOR2X1_430/Y gnd DFFPOSX1_3/D vdd AOI21X1
XDFFPOSX1_19 BUFX2_21/A DFFSR_1/CLK AOI22X1_48/Y gnd vdd DFFPOSX1
XINVX1_157 INVX1_157/A gnd INVX1_157/Y vdd INVX1
XINVX1_146 INVX1_146/A gnd INVX1_146/Y vdd INVX1
XINVX1_168 MUX2X1_29/A gnd INVX1_168/Y vdd INVX1
XINVX1_135 INVX1_135/A gnd INVX1_135/Y vdd INVX1
XINVX1_102 INVX1_102/A gnd INVX1_102/Y vdd INVX1
XINVX1_113 INVX1_113/A gnd INVX1_113/Y vdd INVX1
XINVX1_124 INVX1_124/A gnd INVX1_124/Y vdd INVX1
XINVX1_179 operand_B[45] gnd INVX1_179/Y vdd INVX1
XNOR2X1_504 BUFX4_29/Y AND2X2_74/Y gnd NOR2X1_504/Y vdd NOR2X1
XFILL_32_0_0 gnd vdd FILL
XAOI21X1_117 BUFX4_58/Y INVX1_154/A NOR2X1_185/Y gnd NAND3X1_17/A vdd AOI21X1
XAOI21X1_139 INVX2_75/Y OAI21X1_423/B BUFX4_95/Y gnd OAI21X1_423/C vdd AOI21X1
XAOI21X1_128 BUFX4_186/Y NOR2X1_206/Y NOR2X1_205/Y gnd INVX1_172/A vdd AOI21X1
XAOI21X1_106 BUFX4_184/Y OAI21X1_356/Y NOR2X1_176/Y gnd OR2X2_15/A vdd AOI21X1
XFILL_24_5_1 gnd vdd FILL
XFILL_23_0_0 gnd vdd FILL
XINVX4_10 operand_A[63] gnd INVX4_10/Y vdd INVX4
XINVX4_21 INVX4_21/A gnd INVX4_21/Y vdd INVX4
XFILL_6_1_0 gnd vdd FILL
XFILL_15_5_1 gnd vdd FILL
XFILL_14_0_0 gnd vdd FILL
XNOR2X1_301 NOR2X1_301/A NOR2X1_301/B gnd NOR2X1_301/Y vdd NOR2X1
XNOR2X1_389 NOR2X1_389/A NOR2X1_389/B gnd NOR2X1_389/Y vdd NOR2X1
XFILL_32_1 gnd vdd FILL
XNOR2X1_378 BUFX2_33/A BUFX2_34/A gnd NOR2X1_378/Y vdd NOR2X1
XNOR2X1_312 NOR2X1_312/A NOR2X1_312/B gnd NOR2X1_314/B vdd NOR2X1
XNOR2X1_334 NOR2X1_334/A OAI22X1_17/Y gnd AND2X2_42/A vdd NOR2X1
XNOR2X1_345 INVX2_84/Y INVX2_86/Y gnd NOR2X1_345/Y vdd NOR2X1
XNOR2X1_323 NOR2X1_323/A INVX2_82/Y gnd NOR2X1_323/Y vdd NOR2X1
XNOR2X1_367 OAI22X1_22/D INVX2_91/A gnd INVX1_259/A vdd NOR2X1
XNOR2X1_356 INVX1_255/A INVX1_257/A gnd INVX4_24/A vdd NOR2X1
XOAI21X1_818 OAI21X1_32/A NOR2X1_60/B OAI21X1_30/B gnd NOR2X1_459/B vdd OAI21X1
XOAI21X1_807 OAI21X1_807/A INVX2_17/A BUFX4_140/Y gnd OAI21X1_807/Y vdd OAI21X1
XOAI21X1_829 NOR2X1_462/A NOR2X1_462/B OAI21X1_829/C gnd OAI21X1_829/Y vdd OAI21X1
XNAND3X1_30 NAND3X1_30/A NAND3X1_30/B INVX8_13/Y gnd NAND3X1_30/Y vdd NAND3X1
XNAND3X1_41 NAND3X1_41/A NOR2X1_374/Y NAND3X1_41/C gnd NAND3X1_41/Y vdd NAND3X1
XNOR2X1_30 operand_B[10] INVX2_22/Y gnd NOR2X1_30/Y vdd NOR2X1
XNAND3X1_52 NOR2X1_56/Y AND2X2_46/Y AND2X2_10/Y gnd NOR2X1_413/A vdd NAND3X1
XNAND3X1_63 NAND3X1_63/A NAND3X1_63/B NAND3X1_63/C gnd NOR2X1_454/B vdd NAND3X1
XNOR2X1_96 INVX4_1/Y NOR2X1_96/B gnd NOR2X1_97/B vdd NOR2X1
XNOR2X1_41 INVX4_8/Y INVX1_23/Y gnd NOR2X1_41/Y vdd NOR2X1
XNOR2X1_74 INVX2_34/Y INVX2_36/Y gnd INVX8_7/A vdd NOR2X1
XNOR2X1_85 alu_op[0] INVX2_37/Y gnd INVX1_57/A vdd NOR2X1
XNOR2X1_52 operand_B[20] INVX2_4/Y gnd NOR2X1_52/Y vdd NOR2X1
XNOR2X1_63 operand_B[11] INVX2_27/Y gnd INVX1_83/A vdd NOR2X1
XFILL_30_3_1 gnd vdd FILL
XNAND2X1_7 operand_B[20] INVX2_4/Y gnd NAND2X1_8/B vdd NAND2X1
XNAND2X1_109 BUFX4_20/Y INVX1_46/Y gnd OAI21X1_60/C vdd NAND2X1
XNOR2X1_120 NOR2X1_120/A INVX1_33/Y gnd NOR2X1_120/Y vdd NOR2X1
XMUX2X1_70 operand_A[25] operand_A[24] BUFX4_46/Y gnd MUX2X1_70/Y vdd MUX2X1
XNOR2X1_131 MUX2X1_23/S INVX1_101/Y gnd NAND3X1_7/C vdd NOR2X1
XMUX2X1_81 operand_A[2] operand_A[1] BUFX4_43/Y gnd MUX2X1_83/B vdd MUX2X1
XNOR2X1_142 BUFX4_184/Y INVX1_209/A gnd NOR2X1_142/Y vdd NOR2X1
XNOR2X1_153 operand_A[36] operand_B[36] gnd OAI22X1_5/D vdd NOR2X1
XNOR2X1_164 operand_B[36] INVX2_44/Y gnd NOR2X1_164/Y vdd NOR2X1
XOAI21X1_626 OAI21X1_626/A INVX1_259/Y INVX2_91/Y gnd OAI21X1_626/Y vdd OAI21X1
XOAI21X1_637 OAI22X1_22/D INVX2_91/A INVX4_25/Y gnd OR2X2_38/B vdd OAI21X1
XOAI21X1_604 INVX2_87/Y MUX2X1_7/S OAI21X1_61/C gnd MUX2X1_65/B vdd OAI21X1
XFILL_21_3_1 gnd vdd FILL
XNOR2X1_186 NOR2X1_186/A NOR2X1_186/B gnd AND2X2_15/B vdd NOR2X1
XNOR2X1_175 OR2X2_8/B NOR2X1_175/B gnd NOR2X1_175/Y vdd NOR2X1
XOAI21X1_615 NOR2X1_361/Y NOR2X1_360/Y BUFX4_84/Y gnd NAND3X1_36/C vdd OAI21X1
XNOR2X1_197 BUFX4_41/Y MUX2X1_28/Y gnd NOR2X1_197/Y vdd NOR2X1
XMUX2X1_92 operand_A[10] operand_A[9] BUFX4_50/Y gnd MUX2X1_98/A vdd MUX2X1
XOAI21X1_648 NOR2X1_51/Y NAND2X1_11/B NAND2X1_63/Y gnd OAI21X1_648/Y vdd OAI21X1
XOAI21X1_659 INVX1_204/A OAI21X1_659/B OAI21X1_659/C gnd AOI22X1_30/C vdd OAI21X1
XMUX2X1_126 MUX2X1_126/A MUX2X1_126/B BUFX4_186/Y gnd MUX2X1_126/Y vdd MUX2X1
XMUX2X1_115 MUX2X1_122/B MUX2X1_115/B BUFX4_39/Y gnd MUX2X1_115/Y vdd MUX2X1
XMUX2X1_104 MUX2X1_74/A MUX2X1_71/A MUX2X1_27/S gnd NOR2X1_465/B vdd MUX2X1
XFILL_29_4_1 gnd vdd FILL
XINVX1_77 INVX1_77/A gnd INVX1_77/Y vdd INVX1
XINVX1_22 operand_B[26] gnd INVX1_22/Y vdd INVX1
XINVX1_33 INVX1_33/A gnd INVX1_33/Y vdd INVX1
XNAND2X1_643 BUFX4_184/Y MUX2X1_36/Y gnd OAI21X1_908/C vdd NAND2X1
XINVX1_88 INVX1_88/A gnd INVX1_88/Y vdd INVX1
XINVX1_55 INVX1_55/A gnd INVX1_55/Y vdd INVX1
XNAND2X1_632 operand_B[20] operand_A[20] gnd INVX1_321/A vdd NAND2X1
XINVX1_44 INVX1_44/A gnd INVX1_44/Y vdd INVX1
XFILL_4_4_1 gnd vdd FILL
XINVX1_99 INVX1_99/A gnd INVX1_99/Y vdd INVX1
XINVX1_66 INVX1_66/A gnd INVX1_66/Y vdd INVX1
XNAND2X1_610 OAI21X1_797/Y NOR2X1_453/Y gnd OAI21X1_802/A vdd NAND2X1
XINVX1_11 INVX1_11/A gnd INVX1_11/Y vdd INVX1
XNAND2X1_621 BUFX4_22/Y INVX1_299/A gnd OAI21X1_847/C vdd NAND2X1
XDFFPOSX1_7 BUFX2_9/A CLKBUF1_7/Y DFFPOSX1_7/D gnd vdd DFFPOSX1
XBUFX2_19 BUFX2_19/A gnd result[16] vdd BUFX2
XFILL_12_3_1 gnd vdd FILL
XOAI22X1_17 BUFX4_64/Y INVX1_241/Y BUFX4_157/Y INVX2_84/Y gnd OAI22X1_17/Y vdd OAI22X1
XOAI22X1_28 OAI22X1_28/A OAI22X1_28/B OAI22X1_28/C OAI22X1_28/D gnd AND2X2_68/A vdd
+ OAI22X1
XOAI21X1_478 AND2X2_26/B OAI21X1_565/A OAI21X1_478/C gnd AND2X2_28/B vdd OAI21X1
XOAI21X1_489 OAI21X1_565/A AND2X2_26/B OAI21X1_501/B gnd XNOR2X1_36/A vdd OAI21X1
XOAI21X1_423 INVX2_75/Y OAI21X1_423/B OAI21X1_423/C gnd OAI21X1_423/Y vdd OAI21X1
XOAI21X1_401 BUFX4_75/Y OAI21X1_401/B OAI21X1_401/C gnd MUX2X1_41/B vdd OAI21X1
XOAI21X1_467 INVX1_190/Y MUX2X1_1/S OAI21X1_467/C gnd OAI21X1_467/Y vdd OAI21X1
XOAI21X1_412 INVX2_73/Y BUFX4_43/Y OAI21X1_412/C gnd OAI21X1_412/Y vdd OAI21X1
XOAI21X1_456 INVX2_43/Y BUFX4_48/Y OAI21X1_80/C gnd INVX1_188/A vdd OAI21X1
XOAI21X1_445 operand_A[45] operand_B[45] BUFX4_5/Y gnd NAND3X1_23/A vdd OAI21X1
XOAI21X1_434 INVX1_178/Y NOR2X1_83/A OAI21X1_434/C gnd MUX2X1_47/B vdd OAI21X1
XNAND2X1_462 NOR2X1_265/Y NOR2X1_281/Y gnd NOR2X1_311/B vdd NAND2X1
XNAND2X1_484 AND2X2_35/Y BUFX4_149/Y gnd NAND3X1_33/A vdd NAND2X1
XNAND2X1_451 BUFX4_73/Y INVX1_210/Y gnd OAI21X1_504/C vdd NAND2X1
XNAND2X1_440 MUX2X1_66/S INVX1_217/A gnd OAI21X1_481/C vdd NAND2X1
XNAND2X1_473 BUFX4_19/Y MUX2X1_63/A gnd OAI21X1_537/C vdd NAND2X1
XNAND2X1_495 INVX8_8/A OAI21X1_375/Y gnd OAI21X1_570/C vdd NAND2X1
XFILL_8_2 gnd vdd FILL
XOAI21X1_94 NOR2X1_97/B NOR2X1_97/A OAI21X1_94/C gnd OAI21X1_94/Y vdd OAI21X1
XOAI21X1_61 INVX4_9/Y MUX2X1_1/S OAI21X1_61/C gnd MUX2X1_22/B vdd OAI21X1
XOAI21X1_83 MUX2X1_98/S MUX2X1_9/Y OAI21X1_83/C gnd OAI21X1_83/Y vdd OAI21X1
XOAI21X1_72 INVX1_49/Y BUFX4_68/Y OAI21X1_72/C gnd OAI21X1_72/Y vdd OAI21X1
XOAI21X1_50 BUFX4_17/Y OAI21X1_50/B OAI21X1_50/C gnd OAI22X1_1/C vdd OAI21X1
XFILL_26_2_1 gnd vdd FILL
XFILL_1_2_1 gnd vdd FILL
XOAI21X1_286 INVX4_17/Y OAI22X1_3/D INVX2_62/A gnd INVX1_283/A vdd OAI21X1
XOAI21X1_264 INVX2_60/Y operand_B[34] NAND3X1_9/B gnd XNOR2X1_31/A vdd OAI21X1
XOAI21X1_242 INVX4_15/Y NOR2X1_103/A INVX4_16/A gnd NOR2X1_158/A vdd OAI21X1
XOAI21X1_275 INVX2_61/Y MUX2X1_4/S OAI21X1_275/C gnd OAI21X1_275/Y vdd OAI21X1
XAND2X2_31 AND2X2_31/A INVX8_13/Y gnd AND2X2_31/Y vdd AND2X2
XAND2X2_20 AND2X2_20/A BUFX4_21/Y gnd AND2X2_20/Y vdd AND2X2
XOAI21X1_220 INVX1_106/Y INVX8_3/A OAI21X1_220/C gnd MUX2X1_37/B vdd OAI21X1
XOAI21X1_231 BUFX4_122/Y OAI21X1_231/B OAI21X1_231/C gnd MUX2X1_29/B vdd OAI21X1
XOAI21X1_253 MUX2X1_2/A MUX2X1_2/S OAI21X1_253/C gnd OAI21X1_397/A vdd OAI21X1
XOAI21X1_297 INVX2_58/Y NOR2X1_82/A INVX8_3/A gnd OAI21X1_298/C vdd OAI21X1
XINVX1_306 INVX1_306/A gnd INVX1_306/Y vdd INVX1
XINVX1_328 INVX1_328/A gnd INVX1_328/Y vdd INVX1
XINVX1_317 NOR2X1_10/Y gnd INVX1_317/Y vdd INVX1
XAND2X2_42 AND2X2_42/A INVX8_13/Y gnd AND2X2_42/Y vdd AND2X2
XAND2X2_75 AND2X2_75/A INVX8_7/A gnd AND2X2_75/Y vdd AND2X2
XNAND2X1_270 MUX2X1_99/S OAI21X1_83/Y gnd OAI21X1_246/C vdd NAND2X1
XFILL_9_3_1 gnd vdd FILL
XAND2X2_64 AND2X2_64/A BUFX4_112/Y gnd AND2X2_64/Y vdd AND2X2
XAND2X2_53 AND2X2_53/A AND2X2_53/B gnd AND2X2_53/Y vdd AND2X2
XNAND2X1_281 BUFX4_75/Y OAI21X1_257/Y gnd OAI21X1_258/C vdd NAND2X1
XNAND2X1_292 MUX2X1_51/S INVX1_70/Y gnd OAI21X1_266/C vdd NAND2X1
XFILL_17_2_1 gnd vdd FILL
XINVX1_125 BUFX2_39/A gnd INVX1_125/Y vdd INVX1
XINVX1_169 INVX1_169/A gnd INVX1_169/Y vdd INVX1
XINVX1_158 INVX1_158/A gnd INVX1_158/Y vdd INVX1
XINVX1_103 INVX1_103/A gnd INVX1_103/Y vdd INVX1
XINVX1_136 INVX1_136/A gnd INVX1_136/Y vdd INVX1
XINVX1_114 INVX1_114/A gnd INVX1_114/Y vdd INVX1
XINVX1_147 INVX1_147/A gnd INVX1_147/Y vdd INVX1
XFILL_32_0_1 gnd vdd FILL
XNOR2X1_505 NOR2X1_505/A NOR2X1_505/B gnd NOR2X1_505/Y vdd NOR2X1
XAOI21X1_118 INVX1_154/A INVX1_155/A INVX1_156/A gnd OAI21X1_379/B vdd AOI21X1
XAOI21X1_129 INVX8_18/A INVX1_172/Y OR2X2_20/Y gnd NAND3X1_19/C vdd AOI21X1
XAOI21X1_107 INVX8_2/A AND2X2_7/A NOR2X1_177/Y gnd INVX1_151/A vdd AOI21X1
XFILL_23_0_1 gnd vdd FILL
XINVX4_22 INVX4_22/A gnd INVX4_22/Y vdd INVX4
XINVX4_11 INVX4_11/A gnd INVX4_11/Y vdd INVX4
XFILL_6_1_1 gnd vdd FILL
XFILL_14_0_1 gnd vdd FILL
XNOR2X1_302 BUFX4_98/Y BUFX2_58/A gnd NOR2X1_302/Y vdd NOR2X1
XNOR2X1_313 operand_B[55] INVX2_80/Y gnd NOR2X1_313/Y vdd NOR2X1
XNOR2X1_324 INVX2_81/A INVX2_82/A gnd INVX1_237/A vdd NOR2X1
XNOR2X1_379 BUFX2_35/A BUFX2_36/A gnd NOR2X1_379/Y vdd NOR2X1
XNOR2X1_335 BUFX4_98/Y BUFX2_61/A gnd NOR2X1_335/Y vdd NOR2X1
XNOR2X1_357 INVX1_251/A NOR2X1_357/B gnd NOR2X1_357/Y vdd NOR2X1
XNOR2X1_346 INVX1_198/A OR2X2_17/Y gnd NOR2X1_346/Y vdd NOR2X1
XFILL_25_1 gnd vdd FILL
XNOR2X1_368 OAI22X1_1/B INVX1_261/Y gnd OAI22X1_21/A vdd NOR2X1
XOAI21X1_819 operand_B[10] operand_A[10] BUFX4_1/Y gnd OAI21X1_820/C vdd OAI21X1
XOAI21X1_808 MUX2X1_64/S MUX2X1_127/B NOR2X1_456/Y gnd OAI21X1_810/C vdd OAI21X1
XNAND3X1_42 NOR2X1_381/Y NOR2X1_384/Y NOR2X1_380/Y gnd NOR2X1_394/A vdd NAND3X1
XNAND3X1_31 NAND3X1_31/A NAND3X1_31/B NAND3X1_31/C gnd NAND3X1_31/Y vdd NAND3X1
XNAND3X1_53 NOR2X1_67/Y NAND3X1_53/B NOR2X1_121/Y gnd NAND3X1_54/A vdd NAND3X1
XNOR2X1_42 INVX2_32/Y INVX1_24/Y gnd NOR2X1_42/Y vdd NOR2X1
XNOR2X1_53 operand_B[23] INVX2_8/Y gnd NOR2X1_53/Y vdd NOR2X1
XNAND3X1_20 NAND3X1_20/A NAND3X1_20/B NAND3X1_20/C gnd NAND3X1_20/Y vdd NAND3X1
XNOR2X1_64 operand_B[13] INVX2_20/Y gnd NOR2X1_64/Y vdd NOR2X1
XNOR2X1_20 operand_B[7] INVX1_12/Y gnd INVX1_81/A vdd NOR2X1
XNOR2X1_31 operand_A[10] INVX2_23/Y gnd NOR2X1_31/Y vdd NOR2X1
XNAND3X1_64 XNOR2X1_4/Y INVX1_311/Y INVX1_309/A gnd NAND3X1_65/B vdd NAND3X1
XNOR2X1_97 NOR2X1_97/A NOR2X1_97/B gnd NOR2X1_97/Y vdd NOR2X1
XNOR2X1_86 INVX2_36/Y INVX1_57/Y gnd INVX8_10/A vdd NOR2X1
XNOR2X1_75 NOR2X1_75/A INVX8_7/Y gnd INVX8_8/A vdd NOR2X1
XNAND2X1_8 NAND2X1_8/A NAND2X1_8/B gnd OAI21X1_2/C vdd NAND2X1
XNOR2X1_143 NOR2X1_93/A BUFX2_37/A gnd NOR2X1_143/Y vdd NOR2X1
XNOR2X1_154 OAI22X1_5/D INVX2_63/Y gnd INVX4_19/A vdd NOR2X1
XNOR2X1_121 INVX1_34/A NOR2X1_121/B gnd NOR2X1_121/Y vdd NOR2X1
XNOR2X1_110 NOR2X1_110/A OR2X2_2/Y gnd NOR2X1_110/Y vdd NOR2X1
XMUX2X1_60 MUX2X1_60/A MUX2X1_60/B MUX2X1_62/S gnd MUX2X1_61/B vdd MUX2X1
XMUX2X1_71 MUX2X1_71/A MUX2X1_71/B MUX2X1_71/S gnd MUX2X1_75/B vdd MUX2X1
XNOR2X1_176 BUFX4_183/Y MUX2X1_36/Y gnd NOR2X1_176/Y vdd NOR2X1
XNOR2X1_132 BUFX4_112/Y BUFX4_7/Y gnd INVX4_20/A vdd NOR2X1
XNOR2X1_165 BUFX4_35/Y NOR2X1_165/B gnd INVX1_135/A vdd NOR2X1
XMUX2X1_82 operand_A[4] operand_A[3] MUX2X1_4/S gnd MUX2X1_97/B vdd MUX2X1
XMUX2X1_93 MUX2X1_98/A MUX2X1_93/B BUFX4_66/Y gnd MUX2X1_94/A vdd MUX2X1
XNOR2X1_187 BUFX4_101/Y OR2X2_36/B gnd NOR2X1_187/Y vdd NOR2X1
XOAI21X1_627 OAI21X1_627/A INVX1_259/A NAND3X1_40/B gnd OAI21X1_627/Y vdd OAI21X1
XOAI21X1_616 AND2X2_23/Y INVX2_48/A NOR2X1_80/A gnd OAI21X1_616/Y vdd OAI21X1
XNOR2X1_198 BUFX4_173/Y NOR2X1_198/B gnd NOR2X1_199/B vdd NOR2X1
XOAI21X1_649 OAI21X1_649/A NOR2X1_52/Y NAND2X1_8/B gnd OAI21X1_650/C vdd OAI21X1
XOAI21X1_638 NOR2X1_118/Y NOR2X1_31/Y INVX1_83/Y gnd OAI21X1_640/C vdd OAI21X1
XOAI21X1_605 MUX2X1_32/S INVX1_177/Y OAI21X1_605/C gnd AND2X2_75/A vdd OAI21X1
XMUX2X1_116 MUX2X1_122/A MUX2X1_20/Y BUFX4_21/Y gnd NOR2X1_449/B vdd MUX2X1
XNAND2X1_600 BUFX4_125/Y OAI21X1_708/Y gnd OAI21X1_762/C vdd NAND2X1
XNAND2X1_611 BUFX4_85/Y NOR2X1_195/Y gnd NAND3X1_63/C vdd NAND2X1
XMUX2X1_105 NOR2X1_465/B MUX2X1_121/B BUFX4_24/Y gnd MUX2X1_107/B vdd MUX2X1
XMUX2X1_127 AND2X2_18/A MUX2X1_127/B INVX8_5/A gnd MUX2X1_127/Y vdd MUX2X1
XINVX1_34 INVX1_34/A gnd INVX1_34/Y vdd INVX1
XINVX1_78 INVX1_78/A gnd INVX1_78/Y vdd INVX1
XINVX1_23 operand_B[25] gnd INVX1_23/Y vdd INVX1
XNAND2X1_644 AOI22X1_55/Y OAI22X1_35/Y gnd NAND2X1_644/Y vdd NAND2X1
XINVX1_56 INVX1_56/A gnd INVX1_56/Y vdd INVX1
XNAND2X1_633 INVX2_3/Y INVX2_4/Y gnd AOI22X1_51/D vdd NAND2X1
XINVX1_67 INVX1_67/A gnd INVX1_67/Y vdd INVX1
XINVX1_12 operand_A[7] gnd INVX1_12/Y vdd INVX1
XINVX1_89 INVX1_89/A gnd INVX1_89/Y vdd INVX1
XNAND2X1_622 NAND2X1_622/A AOI22X1_43/Y gnd NAND2X1_622/Y vdd NAND2X1
XINVX1_45 INVX1_45/A gnd INVX1_45/Y vdd INVX1
XDFFPOSX1_8 BUFX2_10/A CLKBUF1_7/Y DFFPOSX1_8/D gnd vdd DFFPOSX1
XAOI21X1_290 NOR2X1_419/Y INVX1_148/A NOR2X1_418/Y gnd OAI21X1_667/C vdd AOI21X1
XOAI22X1_18 INVX2_49/Y OAI22X1_18/B OAI22X1_18/C BUFX4_10/Y gnd OAI22X1_18/Y vdd OAI22X1
XOAI22X1_29 OAI22X1_29/A OAI22X1_29/B OAI22X1_29/C OAI22X1_29/D gnd OAI22X1_29/Y vdd
+ OAI22X1
XOAI21X1_424 OAI21X1_424/A NOR2X1_219/B OAI21X1_424/C gnd OAI21X1_424/Y vdd OAI21X1
XOAI21X1_479 INVX2_42/Y BUFX4_50/Y OAI21X1_71/C gnd OAI21X1_504/B vdd OAI21X1
XOAI21X1_457 BUFX4_73/Y OAI21X1_457/B OAI21X1_457/C gnd MUX2X1_45/B vdd OAI21X1
XOAI21X1_413 INVX1_164/Y BUFX4_69/Y OAI21X1_413/C gnd INVX1_174/A vdd OAI21X1
XOAI21X1_468 INVX1_180/Y BUFX4_69/Y OAI21X1_468/C gnd INVX1_213/A vdd OAI21X1
XOAI21X1_435 BUFX4_163/Y OAI21X1_435/B OAI21X1_435/C gnd OAI21X1_436/C vdd OAI21X1
XOAI21X1_402 MUX2X1_41/B BUFX4_133/Y OAI21X1_402/C gnd MUX2X1_38/B vdd OAI21X1
XOAI21X1_446 INVX1_183/Y BUFX4_39/Y OAI21X1_446/C gnd OAI21X1_945/B vdd OAI21X1
XNAND2X1_463 AND2X2_32/Y BUFX4_153/Y gnd NAND3X1_31/B vdd NAND2X1
XNAND2X1_430 MUX2X1_66/S INVX1_213/A gnd OAI21X1_469/C vdd NAND2X1
XNAND2X1_452 BUFX4_159/Y INVX1_110/A gnd OAI21X1_875/A vdd NAND2X1
XNAND2X1_441 BUFX4_18/Y MUX2X1_54/A gnd OAI21X1_482/C vdd NAND2X1
XNAND2X1_496 BUFX4_116/Y OAI22X1_34/D gnd NAND3X1_34/C vdd NAND2X1
XNAND2X1_485 NAND2X1_485/A OAI21X1_561/Y gnd NAND2X1_485/Y vdd NAND2X1
XNAND2X1_474 INVX2_49/A MUX2X1_34/A gnd OAI21X1_538/C vdd NAND2X1
XOAI21X1_62 MUX2X1_23/S MUX2X1_22/B OAI21X1_62/C gnd OAI21X1_62/Y vdd OAI21X1
XOAI21X1_84 INVX1_50/Y MUX2X1_71/S OAI21X1_84/C gnd OAI21X1_84/Y vdd OAI21X1
XOAI21X1_73 OAI21X1_73/A MUX2X1_30/S OAI21X1_73/C gnd INVX1_146/A vdd OAI21X1
XOAI21X1_51 BUFX4_66/Y INVX2_58/A OAI21X1_51/C gnd MUX2X1_2/B vdd OAI21X1
XOAI21X1_95 INVX4_6/Y BUFX4_50/Y OAI21X1_95/C gnd INVX1_58/A vdd OAI21X1
XOAI21X1_40 INVX4_3/Y MUX2X1_7/S OAI21X1_40/C gnd INVX1_93/A vdd OAI21X1
XOAI21X1_210 INVX1_65/Y BUFX4_74/Y OAI21X1_210/C gnd OAI21X1_315/A vdd OAI21X1
XOAI21X1_221 MUX2X1_34/S MUX2X1_44/B OAI21X1_221/C gnd OAI21X1_222/A vdd OAI21X1
XAND2X2_32 operand_A[52] operand_B[52] gnd AND2X2_32/Y vdd AND2X2
XINVX1_329 NOR2X1_1/Y gnd INVX1_329/Y vdd INVX1
XOAI21X1_243 AOI21X1_62/B NOR2X1_158/A AOI21X1_70/Y gnd OR2X2_9/A vdd OAI21X1
XOAI21X1_287 INVX1_283/A AOI21X1_70/Y AOI21X1_84/Y gnd INVX1_126/A vdd OAI21X1
XAND2X2_43 AND2X2_43/A INVX8_13/Y gnd AND2X2_43/Y vdd AND2X2
XAND2X2_21 operand_A[44] operand_B[44] gnd AND2X2_21/Y vdd AND2X2
XOAI21X1_276 INVX1_105/Y BUFX4_68/Y OAI21X1_276/C gnd INVX1_121/A vdd OAI21X1
XOAI21X1_232 BUFX4_70/Y MUX2X1_13/Y OAI21X1_232/C gnd MUX2X1_28/B vdd OAI21X1
XOAI21X1_265 BUFX4_131/Y OAI21X1_265/B OAI21X1_265/C gnd MUX2X1_39/A vdd OAI21X1
XAND2X2_10 NOR2X1_59/Y NOR2X1_60/Y gnd AND2X2_10/Y vdd AND2X2
XOAI21X1_298 INVX1_90/A NOR2X1_83/A OAI21X1_298/C gnd OR2X2_22/A vdd OAI21X1
XINVX1_307 NOR2X1_35/Y gnd INVX1_307/Y vdd INVX1
XOAI21X1_254 INVX1_45/Y BUFX4_119/Y OAI21X1_254/C gnd INVX1_112/A vdd OAI21X1
XAND2X2_65 AND2X2_65/A AND2X2_65/B gnd AND2X2_65/Y vdd AND2X2
XINVX1_318 INVX1_318/A gnd INVX1_318/Y vdd INVX1
XAND2X2_54 AOI22X1_7/C BUFX4_89/Y gnd AND2X2_54/Y vdd AND2X2
XNAND2X1_293 BUFX4_134/Y INVX1_73/A gnd OAI21X1_268/C vdd NAND2X1
XNAND2X1_271 BUFX4_21/Y MUX2X1_120/B gnd OAI21X1_247/C vdd NAND2X1
XNAND2X1_282 XOR2X1_7/A OAI21X1_48/Y gnd OAI21X1_259/C vdd NAND2X1
XNAND2X1_260 BUFX4_122/Y OAI21X1_308/B gnd OAI21X1_231/C vdd NAND2X1
XFILL_27_5_0 gnd vdd FILL
XFILL_2_5_0 gnd vdd FILL
XFILL_10_4_0 gnd vdd FILL
XINVX1_148 INVX1_148/A gnd INVX1_148/Y vdd INVX1
XINVX1_126 INVX1_126/A gnd INVX1_126/Y vdd INVX1
XINVX1_159 INVX1_159/A gnd INVX1_159/Y vdd INVX1
XINVX1_115 INVX1_115/A gnd INVX1_115/Y vdd INVX1
XINVX1_137 INVX1_137/A gnd INVX1_137/Y vdd INVX1
XINVX1_104 INVX1_104/A gnd INVX1_104/Y vdd INVX1
XNOR2X1_506 NOR2X1_506/A NOR2X1_506/B gnd NOR2X1_506/Y vdd NOR2X1
XFILL_18_5_0 gnd vdd FILL
XAOI21X1_119 INVX1_162/Y OAI21X1_379/B BUFX4_28/Y gnd OAI21X1_379/C vdd AOI21X1
XAOI21X1_108 MUX2X1_57/S INVX1_151/Y NOR2X1_176/Y gnd OR2X2_16/A vdd AOI21X1
XINVX4_23 INVX4_23/A gnd INVX4_23/Y vdd INVX4
XINVX4_12 operand_A[61] gnd INVX4_12/Y vdd INVX4
XNOR2X1_336 BUFX4_98/Y BUFX2_62/A gnd NOR2X1_336/Y vdd NOR2X1
XNOR2X1_303 BUFX4_102/Y BUFX2_59/A gnd NOR2X1_303/Y vdd NOR2X1
XNOR2X1_314 NOR2X1_314/A NOR2X1_314/B gnd INVX1_236/A vdd NOR2X1
XNOR2X1_347 BUFX4_30/Y NOR2X1_357/B gnd NOR2X1_347/Y vdd NOR2X1
XNOR2X1_325 BUFX4_94/Y NOR2X1_325/B gnd NOR2X1_325/Y vdd NOR2X1
XNOR2X1_358 operand_B[60] INVX2_87/Y gnd NOR2X1_359/A vdd NOR2X1
XNOR2X1_369 BUFX4_98/Y BUFX2_65/A gnd NOR2X1_369/Y vdd NOR2X1
XFILL_25_2 gnd vdd FILL
XOAI21X1_809 NOR2X1_196/B BUFX4_77/Y OAI21X1_810/C gnd AOI22X1_38/A vdd OAI21X1
XFILL_24_3_0 gnd vdd FILL
XNAND3X1_21 operand_A[42] INVX2_72/Y NAND3X1_21/C gnd NAND3X1_21/Y vdd NAND3X1
XNAND3X1_32 OR2X2_32/Y NOR2X1_288/Y NAND3X1_32/C gnd NAND3X1_32/Y vdd NAND3X1
XNAND3X1_10 INVX8_13/Y NAND3X1_10/B NAND3X1_10/C gnd NAND3X1_10/Y vdd NAND3X1
XFILL_7_4_0 gnd vdd FILL
XNAND3X1_43 NOR2X1_390/Y NOR2X1_393/Y NOR2X1_389/Y gnd NOR2X1_394/B vdd NAND3X1
XNAND3X1_54 NAND3X1_54/A NAND3X1_54/B NAND3X1_54/C gnd NAND3X1_54/Y vdd NAND3X1
XNOR2X1_43 alu_op[3] alu_op[2] gnd INVX2_33/A vdd NOR2X1
XNOR2X1_87 INVX8_5/A NOR2X1_87/B gnd INVX2_49/A vdd NOR2X1
XNOR2X1_65 operand_B[12] INVX2_21/Y gnd NOR2X1_65/Y vdd NOR2X1
XNOR2X1_32 INVX2_24/Y INVX2_25/Y gnd NOR2X1_32/Y vdd NOR2X1
XNOR2X1_21 operand_A[7] INVX1_13/Y gnd NOR2X1_21/Y vdd NOR2X1
XNOR2X1_76 BUFX4_48/Y INVX1_29/Y gnd INVX2_58/A vdd NOR2X1
XNOR2X1_54 NOR2X1_54/A INVX2_9/Y gnd NOR2X1_54/Y vdd NOR2X1
XNAND3X1_65 BUFX4_105/Y NAND3X1_65/B NAND3X1_65/C gnd NAND3X1_65/Y vdd NAND3X1
XNOR2X1_10 INVX4_5/Y INVX2_5/Y gnd NOR2X1_10/Y vdd NOR2X1
XNOR2X1_98 INVX4_10/Y BUFX4_80/Y gnd INVX1_72/A vdd NOR2X1
XFILL_15_3_0 gnd vdd FILL
XNAND2X1_9 operand_A[18] INVX2_5/Y gnd NAND2X1_9/Y vdd NAND2X1
XNOR2X1_133 NOR2X1_93/A BUFX2_36/A gnd NOR2X1_133/Y vdd NOR2X1
XNOR2X1_144 INVX4_17/Y AND2X2_12/Y gnd NOR2X1_144/Y vdd NOR2X1
XNOR2X1_188 INVX2_54/Y INVX1_161/Y gnd NOR2X1_190/B vdd NOR2X1
XNOR2X1_155 INVX2_62/A OR2X2_9/B gnd NOR2X1_155/Y vdd NOR2X1
XNOR2X1_111 BUFX4_29/Y INVX1_78/Y gnd NOR2X1_111/Y vdd NOR2X1
XMUX2X1_50 MUX2X1_53/B MUX2X1_50/B BUFX4_73/Y gnd MUX2X1_51/B vdd MUX2X1
XNOR2X1_122 INVX1_31/A NOR2X1_122/B gnd NOR2X1_122/Y vdd NOR2X1
XMUX2X1_61 MUX2X1_61/A MUX2X1_61/B INVX8_2/A gnd MUX2X1_61/Y vdd MUX2X1
XNOR2X1_177 BUFX4_42/Y NOR2X1_177/B gnd NOR2X1_177/Y vdd NOR2X1
XNOR2X1_100 MUX2X1_97/S INVX2_57/Y gnd INVX1_73/A vdd NOR2X1
XNOR2X1_199 NOR2X1_199/A NOR2X1_199/B gnd NOR2X1_199/Y vdd NOR2X1
XMUX2X1_83 MUX2X1_97/B MUX2X1_83/B NOR2X1_82/A gnd MUX2X1_87/B vdd MUX2X1
XMUX2X1_94 MUX2X1_94/A MUX2X1_94/B NOR2X1_19/B gnd MUX2X1_95/A vdd MUX2X1
XNOR2X1_166 BUFX4_37/Y NOR2X1_166/B gnd NOR2X1_166/Y vdd NOR2X1
XMUX2X1_72 operand_A[21] operand_A[20] BUFX4_48/Y gnd MUX2X1_72/Y vdd MUX2X1
XOAI21X1_617 BUFX4_157/Y INVX4_24/Y AOI22X1_28/Y gnd NOR2X1_362/B vdd OAI21X1
XOAI21X1_606 OAI21X1_939/A BUFX4_174/Y AND2X2_43/Y gnd OAI21X1_606/Y vdd OAI21X1
XOAI21X1_628 OAI21X1_628/A INVX8_1/A MUX2X1_62/S gnd OAI21X1_628/Y vdd OAI21X1
XOAI21X1_639 INVX1_278/Y NOR2X1_117/Y OAI21X1_639/C gnd OAI21X1_640/A vdd OAI21X1
XINVX1_24 operand_B[24] gnd INVX1_24/Y vdd INVX1
XNAND2X1_645 BUFX4_167/Y NOR2X1_458/B gnd OAI21X1_925/C vdd NAND2X1
XNAND2X1_634 OAI21X1_886/Y NOR2X1_492/Y gnd NAND2X1_634/Y vdd NAND2X1
XMUX2X1_128 MUX2X1_39/Y NOR2X1_461/B OR2X2_43/B gnd MUX2X1_128/Y vdd MUX2X1
XNAND2X1_623 BUFX4_184/Y OAI21X1_86/B gnd NAND2X1_623/Y vdd NAND2X1
XMUX2X1_117 MUX2X1_24/Y MUX2X1_75/B BUFX4_42/Y gnd MUX2X1_126/B vdd MUX2X1
XINVX1_13 operand_B[7] gnd INVX1_13/Y vdd INVX1
XMUX2X1_106 MUX2X1_106/A MUX2X1_74/B BUFX4_125/Y gnd NOR2X1_464/B vdd MUX2X1
XNAND2X1_612 XOR2X1_4/A OAI21X1_727/A gnd OAI21X1_814/C vdd NAND2X1
XNAND2X1_601 OR2X2_39/B NOR2X1_471/B gnd OAI21X1_763/C vdd NAND2X1
XINVX1_35 alu_op[0] gnd INVX1_35/Y vdd INVX1
XINVX1_57 INVX1_57/A gnd INVX1_57/Y vdd INVX1
XINVX1_68 INVX1_68/A gnd INVX1_68/Y vdd INVX1
XINVX1_79 MUX2X1_7/S gnd INVX1_79/Y vdd INVX1
XINVX1_46 INVX1_46/A gnd INVX1_46/Y vdd INVX1
XDFFPOSX1_9 BUFX2_11/A CLKBUF1_2/Y DFFPOSX1_9/D gnd vdd DFFPOSX1
XAOI21X1_291 INVX1_283/Y OAI21X1_666/Y OAI21X1_665/Y gnd NOR2X1_420/B vdd AOI21X1
XAOI21X1_280 INVX1_30/A INVX2_19/Y INVX1_85/Y gnd AND2X2_48/B vdd AOI21X1
XFILL_30_1_0 gnd vdd FILL
XFILL_21_1_0 gnd vdd FILL
XOAI21X1_414 INVX1_174/Y MUX2X1_87/S OAI21X1_414/C gnd INVX1_175/A vdd OAI21X1
XOAI21X1_403 MUX2X1_57/A BUFX4_183/Y BUFX4_79/Y gnd OAI21X1_404/B vdd OAI21X1
XOAI22X1_19 OAI22X1_19/A OAI22X1_1/B OAI22X1_19/C INVX8_8/Y gnd OAI22X1_37/D vdd OAI22X1
XOAI21X1_425 NOR2X1_217/A AND2X2_21/Y NOR2X1_220/B gnd OAI21X1_425/Y vdd OAI21X1
XOAI21X1_436 NOR2X1_467/B OR2X2_25/B OAI21X1_436/C gnd OR2X2_23/B vdd OAI21X1
XOAI21X1_469 INVX1_174/Y BUFX4_120/Y OAI21X1_469/C gnd OAI21X1_469/Y vdd OAI21X1
XOAI21X1_447 AND2X2_23/Y INVX2_48/A BUFX4_184/Y gnd OAI21X1_448/C vdd OAI21X1
XOAI21X1_458 INVX1_187/Y BUFX4_19/Y OAI21X1_458/C gnd INVX1_261/A vdd OAI21X1
XNAND2X1_486 INVX2_79/A INVX1_224/A gnd NOR2X1_307/A vdd NAND2X1
XNAND2X1_475 INVX2_78/A INVX1_219/A gnd NOR2X1_307/B vdd NAND2X1
XNAND2X1_453 operand_A[50] INVX2_76/Y gnd OAI21X1_520/B vdd NAND2X1
XNAND2X1_464 BUFX4_159/Y INVX1_133/A gnd OAI22X1_12/B vdd NAND2X1
XNAND2X1_497 NOR2X1_80/A OAI21X1_391/Y gnd NAND2X1_497/Y vdd NAND2X1
XNAND2X1_431 BUFX4_19/Y OAI21X1_469/Y gnd OAI21X1_470/C vdd NAND2X1
XNAND2X1_442 BUFX4_164/Y INVX1_86/A gnd NOR2X1_252/B vdd NAND2X1
XNAND2X1_420 BUFX4_186/Y NOR2X1_228/Y gnd OAI21X1_449/C vdd NAND2X1
XFILL_29_2_0 gnd vdd FILL
XFILL_4_2_0 gnd vdd FILL
XFILL_12_1_0 gnd vdd FILL
XOAI21X1_63 INVX2_38/Y MUX2X1_6/S OAI21X1_63/C gnd INVX1_47/A vdd OAI21X1
XOAI21X1_52 INVX4_7/Y MUX2X1_6/S OAI21X1_52/C gnd OAI21X1_54/B vdd OAI21X1
XOAI21X1_30 NOR2X1_60/A OAI21X1_30/B OAI21X1_30/C gnd OAI21X1_30/Y vdd OAI21X1
XOAI21X1_41 INVX1_38/Y BUFX4_67/Y OAI21X1_41/C gnd INVX1_113/A vdd OAI21X1
XOAI21X1_74 BUFX4_39/Y INVX1_146/A OAI21X1_74/C gnd OAI21X1_74/Y vdd OAI21X1
XOAI21X1_85 BUFX4_41/Y OAI21X1_85/B OAI21X1_85/C gnd OAI21X1_86/B vdd OAI21X1
XOAI21X1_96 INVX2_7/Y MUX2X1_7/S OAI21X1_96/C gnd OAI21X1_96/Y vdd OAI21X1
XOAI21X1_244 INVX4_17/Y OAI22X1_3/D OR2X2_9/A gnd NAND3X1_9/B vdd OAI21X1
XOAI21X1_200 INVX1_96/Y BUFX4_120/Y OAI21X1_200/C gnd OAI21X1_374/B vdd OAI21X1
XOAI21X1_233 INVX2_57/Y BUFX4_67/Y OAI21X1_312/A gnd MUX2X1_28/A vdd OAI21X1
XOAI21X1_211 BUFX4_190/Y OAI21X1_211/B OAI21X1_211/C gnd MUX2X1_35/B vdd OAI21X1
XOAI21X1_255 BUFX4_20/Y OAI21X1_397/A OAI21X1_255/C gnd OAI21X1_261/B vdd OAI21X1
XOAI21X1_222 OAI21X1_222/A BUFX4_111/Y OAI21X1_222/C gnd NAND3X1_8/C vdd OAI21X1
XAND2X2_33 operand_A[54] operand_B[54] gnd AND2X2_33/Y vdd AND2X2
XAND2X2_44 operand_A[63] operand_B[63] gnd AND2X2_44/Y vdd AND2X2
XOAI21X1_288 AOI21X1_62/B INVX1_127/Y INVX1_126/Y gnd INVX1_144/A vdd OAI21X1
XOAI21X1_266 BUFX4_133/Y MUX2X1_20/B OAI21X1_266/C gnd INVX1_117/A vdd OAI21X1
XAND2X2_55 AND2X2_55/A INVX8_12/A gnd AND2X2_55/Y vdd AND2X2
XOAI21X1_299 BUFX4_131/Y OAI21X1_299/B OAI21X1_299/C gnd MUX2X1_33/A vdd OAI21X1
XAND2X2_22 AND2X2_22/A BUFX4_159/Y gnd OR2X2_44/A vdd AND2X2
XINVX1_308 BUFX2_15/A gnd INVX1_308/Y vdd INVX1
XAND2X2_66 AND2X2_66/A AND2X2_66/B gnd AND2X2_66/Y vdd AND2X2
XAND2X2_11 AND2X2_11/A AND2X2_11/B gnd OR2X2_5/A vdd AND2X2
XINVX1_319 NOR2X1_9/Y gnd INVX1_319/Y vdd INVX1
XOAI21X1_277 INVX1_121/Y BUFX4_131/Y OAI21X1_277/C gnd OAI21X1_415/B vdd OAI21X1
XNAND2X1_250 INVX8_1/A OAI21X1_103/Y gnd OAI21X1_219/C vdd NAND2X1
XNAND2X1_294 BUFX4_38/Y OAI21X1_268/Y gnd OAI21X1_269/C vdd NAND2X1
XNAND2X1_272 BUFX4_159/Y MUX2X1_124/B gnd AOI21X1_72/A vdd NAND2X1
XNAND2X1_261 BUFX4_22/Y MUX2X1_29/B gnd OAI21X1_234/C vdd NAND2X1
XNAND2X1_283 BUFX4_18/Y MUX2X1_38/A gnd OAI21X1_260/C vdd NAND2X1
XFILL_6_1 gnd vdd FILL
XFILL_27_5_1 gnd vdd FILL
XFILL_26_0_0 gnd vdd FILL
XFILL_2_5_1 gnd vdd FILL
XFILL_1_0_0 gnd vdd FILL
XINVX1_116 operand_B[35] gnd INVX1_116/Y vdd INVX1
XINVX1_105 INVX1_105/A gnd INVX1_105/Y vdd INVX1
XFILL_10_4_1 gnd vdd FILL
XINVX1_127 INVX1_127/A gnd INVX1_127/Y vdd INVX1
XINVX1_149 INVX1_149/A gnd INVX1_149/Y vdd INVX1
XINVX1_138 INVX1_138/A gnd INVX1_138/Y vdd INVX1
XFILL_9_1_0 gnd vdd FILL
XNOR2X1_507 NOR2X1_93/A BUFX2_31/A gnd NOR2X1_507/Y vdd NOR2X1
XFILL_18_5_1 gnd vdd FILL
XFILL_17_0_0 gnd vdd FILL
XAOI21X1_109 INVX8_11/A XNOR2X1_33/Y NAND3X1_15/Y gnd AOI21X1_110/A vdd AOI21X1
XINVX4_24 INVX4_24/A gnd INVX4_24/Y vdd INVX4
XINVX4_13 operand_A[57] gnd INVX4_13/Y vdd INVX4
XNOR2X1_326 BUFX4_98/Y OR2X2_37/B gnd NOR2X1_326/Y vdd NOR2X1
XNOR2X1_348 INVX2_84/A OR2X2_34/B gnd INVX1_249/A vdd NOR2X1
XNOR2X1_337 INVX2_85/Y INVX1_242/Y gnd INVX1_243/A vdd NOR2X1
XNOR2X1_304 operand_A[56] operand_B[56] gnd NOR2X1_306/A vdd NOR2X1
XNOR2X1_359 NOR2X1_359/A INVX4_24/Y gnd NOR2X1_359/Y vdd NOR2X1
XNOR2X1_315 NOR2X1_75/A MUX2X1_54/Y gnd NOR2X1_315/Y vdd NOR2X1
XFILL_24_3_1 gnd vdd FILL
XNAND3X1_33 NAND3X1_33/A NAND3X1_33/B INVX8_13/Y gnd NAND3X1_33/Y vdd NAND3X1
XNAND3X1_11 AOI22X1_4/C INVX4_16/Y NOR2X1_155/Y gnd OR2X2_17/A vdd NAND3X1
XNAND3X1_55 INVX2_90/Y operand_B[62] INVX4_25/Y gnd AND2X2_50/A vdd NAND3X1
XNAND3X1_22 NAND3X1_22/A NOR2X1_224/Y NAND3X1_22/C gnd OR2X2_23/A vdd NAND3X1
XNAND3X1_44 INVX1_262/Y INVX1_263/Y NOR2X1_395/Y gnd NOR2X1_397/A vdd NAND3X1
XFILL_7_4_1 gnd vdd FILL
XNAND3X1_66 NAND3X1_66/A NAND3X1_66/B NAND3X1_66/C gnd NAND3X1_66/Y vdd NAND3X1
XNOR2X1_44 alu_op[1] alu_op[0] gnd INVX1_27/A vdd NOR2X1
XNOR2X1_99 MUX2X1_6/S INVX4_10/Y gnd INVX2_57/A vdd NOR2X1
XNOR2X1_11 INVX2_8/Y INVX1_8/Y gnd NOR2X1_11/Y vdd NOR2X1
XNOR2X1_88 INVX2_33/Y INVX1_51/Y gnd BUFX4_6/A vdd NOR2X1
XNOR2X1_77 INVX2_37/Y INVX2_36/Y gnd INVX8_9/A vdd NOR2X1
XFILL_15_3_1 gnd vdd FILL
XNOR2X1_33 INVX2_26/Y INVX1_20/Y gnd NOR2X1_33/Y vdd NOR2X1
XNOR2X1_55 BUFX4_36/Y INVX2_11/Y gnd INVX1_80/A vdd NOR2X1
XNOR2X1_22 NOR2X1_22/A INVX2_14/Y gnd NOR2X1_22/Y vdd NOR2X1
XNOR2X1_66 NOR2X1_66/A NOR2X1_66/B gnd NOR2X1_66/Y vdd NOR2X1
XFILL_30_1 gnd vdd FILL
XNOR2X1_123 operand_B[31] INVX2_50/Y gnd NOR2X1_123/Y vdd NOR2X1
XNOR2X1_134 operand_A[34] operand_B[34] gnd OAI22X1_3/D vdd NOR2X1
XNOR2X1_156 operand_B[34] INVX2_60/Y gnd NOR2X1_156/Y vdd NOR2X1
XNOR2X1_178 INVX2_47/Y INVX1_152/Y gnd INVX1_156/A vdd NOR2X1
XNOR2X1_189 operand_A[41] operand_B[41] gnd NOR2X1_190/A vdd NOR2X1
XNOR2X1_167 OR2X2_8/B NOR2X1_167/B gnd NOR2X1_167/Y vdd NOR2X1
XMUX2X1_51 MUX2X1_51/A MUX2X1_51/B MUX2X1_51/S gnd MUX2X1_67/A vdd MUX2X1
XMUX2X1_62 MUX2X1_62/A MUX2X1_62/B MUX2X1_62/S gnd MUX2X1_63/B vdd MUX2X1
XMUX2X1_73 operand_A[23] operand_A[22] MUX2X1_1/S gnd MUX2X1_73/Y vdd MUX2X1
XNOR2X1_101 BUFX4_136/Y INVX1_73/Y gnd AND2X2_7/A vdd NOR2X1
XMUX2X1_40 MUX2X1_47/B MUX2X1_40/B BUFX4_18/Y gnd MUX2X1_40/Y vdd MUX2X1
XMUX2X1_84 operand_A[8] operand_A[7] MUX2X1_9/S gnd MUX2X1_98/B vdd MUX2X1
XNOR2X1_112 operand_A[0] INVX1_79/Y gnd NOR2X1_112/Y vdd NOR2X1
XMUX2X1_95 MUX2X1_95/A MUX2X1_95/B BUFX4_39/Y gnd MUX2X1_95/Y vdd MUX2X1
XNOR2X1_145 MUX2X1_57/S NOR2X1_145/B gnd NOR2X1_145/Y vdd NOR2X1
XOAI21X1_618 OAI21X1_946/A BUFX4_174/Y NOR2X1_362/Y gnd OAI21X1_618/Y vdd OAI21X1
XOAI21X1_607 OAI21X1_607/A OR2X2_40/B OAI21X1_607/C gnd NOR2X1_352/A vdd OAI21X1
XOAI21X1_629 NOR2X1_54/A INVX2_57/Y OAI21X1_629/C gnd OAI21X1_630/C vdd OAI21X1
XMUX2X1_129 AND2X2_22/A MUX2X1_129/B BUFX4_179/Y gnd MUX2X1_129/Y vdd MUX2X1
XMUX2X1_118 MUX2X1_118/A MUX2X1_27/Y BUFX4_24/Y gnd MUX2X1_127/B vdd MUX2X1
XMUX2X1_107 MUX2X1_107/A MUX2X1_107/B MUX2X1_25/S gnd MUX2X1_107/Y vdd MUX2X1
XINVX1_25 INVX1_25/A gnd INVX1_25/Y vdd INVX1
XNAND2X1_646 NOR2X1_500/Y OAI22X1_36/Y gnd NOR2X1_501/B vdd NAND2X1
XINVX1_47 INVX1_47/A gnd INVX1_47/Y vdd INVX1
XNAND2X1_635 BUFX2_23/A BUFX4_12/Y gnd OAI21X1_890/C vdd NAND2X1
XINVX1_14 operand_B[6] gnd INVX1_14/Y vdd INVX1
XINVX1_36 INVX1_36/A gnd INVX1_36/Y vdd INVX1
XINVX1_58 INVX1_58/A gnd INVX1_58/Y vdd INVX1
XNAND2X1_602 BUFX4_125/Y INVX1_291/A gnd OAI21X1_768/C vdd NAND2X1
XNAND2X1_613 XNOR2X1_7/Y NOR2X1_459/B gnd OAI21X1_824/C vdd NAND2X1
XNAND2X1_624 operand_B[14] operand_A[14] gnd OAI21X1_855/B vdd NAND2X1
XINVX1_69 INVX1_69/A gnd INVX1_69/Y vdd INVX1
XAOI21X1_270 INVX4_20/A AND2X2_3/A NAND2X1_523/Y gnd NAND2X1_524/A vdd AOI21X1
XAOI21X1_292 OAI21X1_671/Y NAND2X1_555/Y OR2X2_29/A gnd NOR2X1_423/B vdd AOI21X1
XAOI21X1_281 AOI22X1_29/Y AND2X2_48/Y OAI21X1_168/B gnd OAI21X1_655/B vdd AOI21X1
XFILL_30_1_1 gnd vdd FILL
XFILL_21_1_1 gnd vdd FILL
XOAI21X1_437 INVX4_21/A NOR2X1_226/Y OAI21X1_437/C gnd OAI21X1_437/Y vdd OAI21X1
XOAI21X1_426 MUX2X1_33/A OR2X2_13/B OAI21X1_426/C gnd AND2X2_22/A vdd OAI21X1
XOAI21X1_448 OAI21X1_945/B MUX2X1_57/S OAI21X1_448/C gnd AND2X2_63/A vdd OAI21X1
XOAI21X1_404 NOR2X1_204/Y OAI21X1_404/B OAI21X1_404/C gnd NAND3X1_19/A vdd OAI21X1
XOAI21X1_415 BUFX4_19/Y OAI21X1_415/B OAI21X1_415/C gnd NOR2X1_212/B vdd OAI21X1
XOAI21X1_459 OAI22X1_1/C MUX2X1_32/S OAI21X1_459/C gnd OAI21X1_460/A vdd OAI21X1
XNAND2X1_487 NOR2X1_307/Y NOR2X1_278/Y gnd INVX1_231/A vdd NAND2X1
XNAND2X1_476 INVX1_224/A INVX1_225/A gnd NAND2X1_476/Y vdd NAND2X1
XFILL_29_2_1 gnd vdd FILL
XNAND2X1_443 operand_A[48] INVX1_197/Y gnd OAI21X1_501/B vdd NAND2X1
XNAND2X1_410 INVX2_75/Y OAI21X1_423/B gnd OAI21X1_454/A vdd NAND2X1
XNAND2X1_432 INVX1_186/A INVX4_22/Y gnd OR2X2_28/A vdd NAND2X1
XNAND2X1_421 INVX2_75/A INVX4_21/Y gnd NOR2X1_244/A vdd NAND2X1
XNAND2X1_454 BUFX4_69/Y OAI21X1_511/Y gnd OAI21X1_512/C vdd NAND2X1
XNAND2X1_498 BUFX4_184/Y MUX2X1_37/Y gnd NAND2X1_498/Y vdd NAND2X1
XFILL_4_2_1 gnd vdd FILL
XNAND2X1_465 MUX2X1_32/S MUX2X1_32/B gnd OAI21X1_524/C vdd NAND2X1
XFILL_12_1_1 gnd vdd FILL
XINVX2_90 operand_A[62] gnd INVX2_90/Y vdd INVX2
XOAI21X1_75 INVX2_44/Y BUFX4_50/Y OAI21X1_75/C gnd OAI21X1_76/B vdd OAI21X1
XOAI21X1_64 INVX2_39/Y BUFX4_53/Y OAI21X1_64/C gnd MUX2X1_22/A vdd OAI21X1
XOAI21X1_20 INVX2_29/Y INVX2_30/Y OAI21X1_20/C gnd OAI21X1_21/C vdd OAI21X1
XOAI21X1_86 MUX2X1_57/S OAI21X1_86/B OAI21X1_86/C gnd OAI21X1_86/Y vdd OAI21X1
XOAI21X1_31 NOR2X1_59/A INVX1_84/A OAI21X1_31/C gnd OAI21X1_31/Y vdd OAI21X1
XOAI21X1_53 INVX2_13/Y BUFX4_53/Y OAI21X1_53/C gnd INVX1_44/A vdd OAI21X1
XOAI21X1_42 INVX1_37/Y BUFX4_119/Y OAI21X1_42/C gnd OAI21X1_50/B vdd OAI21X1
XOAI21X1_97 INVX1_58/Y BUFX4_76/Y OAI21X1_97/C gnd INVX1_59/A vdd OAI21X1
XOAI21X1_289 INVX4_19/Y INVX1_144/A AOI21X1_85/Y gnd OAI21X1_289/Y vdd OAI21X1
XOAI21X1_223 BUFX4_190/Y OAI21X1_223/B OAI21X1_223/C gnd OAI21X1_225/B vdd OAI21X1
XOAI21X1_245 MUX2X1_30/S OAI21X1_72/Y OAI21X1_245/C gnd OAI21X1_247/A vdd OAI21X1
XOAI21X1_234 BUFX4_22/Y MUX2X1_28/Y OAI21X1_234/C gnd OAI21X1_234/Y vdd OAI21X1
XOAI21X1_212 BUFX4_125/Y OAI21X1_315/A OAI21X1_212/C gnd INVX1_103/A vdd OAI21X1
XOAI21X1_256 INVX1_113/Y BUFX4_119/Y OAI21X1_256/C gnd INVX1_114/A vdd OAI21X1
XOAI21X1_278 INVX1_120/Y BUFX4_19/Y OAI21X1_278/C gnd MUX2X1_46/B vdd OAI21X1
XOAI21X1_201 INVX1_94/Y BUFX4_17/Y OAI21X1_201/C gnd MUX2X1_42/B vdd OAI21X1
XOAI21X1_267 INVX1_117/Y BUFX4_37/Y OAI21X1_267/C gnd NOR2X1_145/B vdd OAI21X1
XAND2X2_45 AND2X2_45/A AND2X2_45/B gnd BUFX2_67/A vdd AND2X2
XAND2X2_12 AND2X2_12/A INVX2_59/A gnd AND2X2_12/Y vdd AND2X2
XAND2X2_34 AND2X2_34/A INVX8_13/Y gnd AND2X2_34/Y vdd AND2X2
XAND2X2_23 AND2X2_23/A BUFX4_21/Y gnd AND2X2_23/Y vdd AND2X2
XINVX1_309 INVX1_309/A gnd INVX1_309/Y vdd INVX1
XAND2X2_67 AND2X2_67/A AND2X2_67/B gnd AND2X2_67/Y vdd AND2X2
XAND2X2_56 AND2X2_56/A BUFX4_116/Y gnd AND2X2_56/Y vdd AND2X2
XNAND2X1_262 BUFX4_70/Y OAI21X1_126/Y gnd OAI21X1_232/C vdd NAND2X1
XNAND2X1_273 MUX2X1_51/S OAI21X1_66/B gnd OAI21X1_248/C vdd NAND2X1
XNAND2X1_251 XOR2X1_7/A OAI21X1_219/Y gnd OAI21X1_220/C vdd NAND2X1
XNAND2X1_240 BUFX4_76/Y INVX1_58/A gnd OAI21X1_208/C vdd NAND2X1
XNAND2X1_295 BUFX4_24/Y NOR2X1_147/Y gnd OR2X2_10/A vdd NAND2X1
XNAND2X1_284 MUX2X1_25/S OAI21X1_506/A gnd OAI21X1_261/C vdd NAND2X1
XOAI21X1_790 INVX8_15/Y NAND3X1_14/Y OAI21X1_790/C gnd NOR2X1_451/B vdd OAI21X1
XFILL_26_0_1 gnd vdd FILL
XFILL_1_0_1 gnd vdd FILL
XINVX1_106 INVX1_106/A gnd INVX1_106/Y vdd INVX1
XINVX1_139 INVX1_139/A gnd INVX1_139/Y vdd INVX1
XINVX1_128 INVX1_128/A gnd INVX1_128/Y vdd INVX1
XINVX1_117 INVX1_117/A gnd INVX1_117/Y vdd INVX1
XFILL_9_1_1 gnd vdd FILL
XNOR2X1_508 NOR2X1_2/Y AND2X2_74/Y gnd NOR2X1_508/Y vdd NOR2X1
XFILL_17_0_1 gnd vdd FILL
XINVX4_25 INVX4_25/A gnd INVX4_25/Y vdd INVX4
XINVX4_14 operand_A[45] gnd INVX4_14/Y vdd INVX4
XNOR2X1_327 operand_A[58] operand_B[58] gnd NOR2X1_333/A vdd NOR2X1
XNOR2X1_338 operand_A[59] operand_B[59] gnd INVX1_244/A vdd NOR2X1
XNOR2X1_349 operand_B[59] INVX2_85/Y gnd NOR2X1_349/Y vdd NOR2X1
XNOR2X1_305 INVX2_39/Y INVX1_230/Y gnd NOR2X1_321/A vdd NOR2X1
XNOR2X1_316 BUFX4_167/Y NOR2X1_316/B gnd NOR2X1_316/Y vdd NOR2X1
XNAND3X1_23 NAND3X1_23/A NAND3X1_23/B INVX8_13/Y gnd NAND3X1_23/Y vdd NAND3X1
XNAND3X1_12 NAND3X1_12/A NAND3X1_12/B NAND3X1_12/C gnd NOR2X1_162/B vdd NAND3X1
XNAND3X1_34 INVX8_13/Y AND2X2_37/Y NAND3X1_34/C gnd NAND3X1_34/Y vdd NAND3X1
XNOR2X1_12 INVX1_9/Y INVX4_3/Y gnd OR2X2_49/B vdd NOR2X1
XNAND3X1_67 BUFX4_138/Y NAND3X1_67/B OR2X2_45/Y gnd NAND3X1_68/A vdd NAND3X1
XNAND3X1_56 MUX2X1_64/S NAND3X1_56/B NAND3X1_56/C gnd NAND3X1_56/Y vdd NAND3X1
XNAND3X1_45 INVX1_264/Y INVX1_265/Y NOR2X1_396/Y gnd NOR2X1_397/B vdd NAND3X1
XNOR2X1_67 NOR2X1_67/A NOR2X1_67/B gnd NOR2X1_67/Y vdd NOR2X1
XNOR2X1_45 INVX2_33/Y INVX1_27/Y gnd NOR2X1_45/Y vdd NOR2X1
XNOR2X1_78 INVX2_37/Y INVX1_35/Y gnd INVX1_51/A vdd NOR2X1
XNOR2X1_89 INVX2_33/Y INVX1_57/Y gnd NOR2X1_89/Y vdd NOR2X1
XNOR2X1_56 OR2X2_3/A OR2X2_3/B gnd NOR2X1_56/Y vdd NOR2X1
XNOR2X1_34 INVX2_27/Y INVX2_28/Y gnd NOR2X1_34/Y vdd NOR2X1
XNOR2X1_23 operand_A[5] BUFX4_82/Y gnd NOR2X1_23/Y vdd NOR2X1
XNOR2X1_102 operand_A[32] operand_B[32] gnd NOR2X1_103/A vdd NOR2X1
XMUX2X1_30 MUX2X1_30/A MUX2X1_30/B MUX2X1_30/S gnd MUX2X1_39/B vdd MUX2X1
XMUX2X1_41 MUX2X1_45/B MUX2X1_41/B MUX2X1_66/S gnd MUX2X1_52/A vdd MUX2X1
XMUX2X1_63 MUX2X1_63/A MUX2X1_63/B XOR2X1_4/A gnd MUX2X1_63/Y vdd MUX2X1
XMUX2X1_52 MUX2X1_52/A MUX2X1_67/A XOR2X1_4/A gnd MUX2X1_52/Y vdd MUX2X1
XNOR2X1_113 XOR2X1_7/Y XOR2X1_4/Y gnd AND2X2_46/B vdd NOR2X1
XNOR2X1_124 NOR2X1_22/A INVX8_9/Y gnd AND2X2_11/B vdd NOR2X1
XOAI21X1_608 INVX4_24/Y NOR2X1_357/Y OAI21X1_608/C gnd OAI21X1_608/Y vdd OAI21X1
XFILL_30_2 gnd vdd FILL
XNOR2X1_135 OAI22X1_3/D INVX4_17/Y gnd INVX2_59/A vdd NOR2X1
XNOR2X1_157 operand_B[35] INVX2_61/Y gnd NOR2X1_157/Y vdd NOR2X1
XOAI21X1_619 INVX1_251/Y INVX1_255/A INVX1_257/Y gnd OAI21X1_621/B vdd OAI21X1
XNOR2X1_179 operand_A[40] operand_B[40] gnd NOR2X1_185/A vdd NOR2X1
XFILL_23_1 gnd vdd FILL
XNOR2X1_146 BUFX4_173/Y NOR2X1_435/B gnd NOR2X1_149/B vdd NOR2X1
XMUX2X1_85 operand_A[6] operand_A[5] BUFX4_46/Y gnd MUX2X1_97/A vdd MUX2X1
XMUX2X1_96 MUX2X1_96/A MUX2X1_96/B OR2X2_13/B gnd MUX2X1_96/Y vdd MUX2X1
XMUX2X1_74 MUX2X1_74/A MUX2X1_74/B INVX8_3/A gnd MUX2X1_75/A vdd MUX2X1
XNOR2X1_168 BUFX4_173/Y MUX2X1_34/Y gnd NOR2X1_168/Y vdd NOR2X1
XMUX2X1_108 MUX2X1_94/A MUX2X1_87/A MUX2X1_87/S gnd MUX2X1_109/B vdd MUX2X1
XMUX2X1_119 MUX2X1_119/A MUX2X1_95/A INVX8_2/A gnd NOR2X1_455/B vdd MUX2X1
XINVX1_26 INVX1_26/A gnd INVX1_26/Y vdd INVX1
XNAND2X1_647 XNOR2X1_27/Y OAI21X1_924/A gnd OAI21X1_932/C vdd NAND2X1
XINVX1_48 INVX1_48/A gnd INVX1_48/Y vdd INVX1
XINVX1_15 operand_B[15] gnd INVX1_15/Y vdd INVX1
XINVX1_59 INVX1_59/A gnd INVX1_59/Y vdd INVX1
XNAND2X1_614 BUFX4_138/Y OAI21X1_824/C gnd OAI21X1_822/A vdd NAND2X1
XNAND2X1_603 BUFX4_37/Y OAI21X1_852/B gnd OAI21X1_769/C vdd NAND2X1
XNAND2X1_625 BUFX2_17/A BUFX4_11/Y gnd OAI21X1_856/C vdd NAND2X1
XINVX1_37 INVX1_37/A gnd INVX1_37/Y vdd INVX1
XNAND2X1_636 BUFX4_162/Y NOR2X1_442/B gnd OAI21X1_894/C vdd NAND2X1
XAOI21X1_271 AOI21X1_271/A NAND3X1_40/C NAND2X1_524/Y gnd AOI21X1_272/B vdd AOI21X1
XAOI21X1_293 INVX1_200/A OAI21X1_667/Y OAI21X1_673/Y gnd OAI21X1_674/A vdd AOI21X1
XAOI21X1_260 INVX4_11/Y OAI21X1_616/Y BUFX4_8/Y gnd NOR2X1_509/A vdd AOI21X1
XAOI21X1_282 OAI21X1_647/Y INVX1_282/Y OAI21X1_648/Y gnd OAI21X1_649/A vdd AOI21X1
XOAI21X1_438 INVX2_46/Y operand_B[44] OAI21X1_454/A gnd XNOR2X1_34/A vdd OAI21X1
XOAI21X1_427 XOR2X1_7/A BUFX4_42/Y operand_A[63] gnd INVX1_250/A vdd OAI21X1
XOAI21X1_405 BUFX4_16/Y OAI21X1_405/B OAI21X1_405/C gnd INVX1_324/A vdd OAI21X1
XOAI21X1_449 OAI21X1_945/B INVX8_5/A OAI21X1_449/C gnd AND2X2_64/A vdd OAI21X1
XOAI21X1_416 NOR2X1_211/Y NOR2X1_212/Y BUFX4_84/Y gnd NAND3X1_20/B vdd OAI21X1
XNAND2X1_400 INVX1_169/A INVX2_74/A gnd NOR2X1_219/B vdd NAND2X1
XNAND2X1_411 XOR2X1_4/A INVX1_137/Y gnd OAI21X1_439/C vdd NAND2X1
XNAND2X1_488 NOR2X1_307/Y OAI21X1_518/Y gnd AND2X2_36/A vdd NAND2X1
XNAND2X1_433 NOR2X1_219/Y NOR2X1_244/Y gnd INVX1_198/A vdd NAND2X1
XNAND2X1_444 MUX2X1_6/S operand_A[48] gnd OAI21X1_491/C vdd NAND2X1
XNAND2X1_466 BUFX4_73/Y MUX2X1_50/B gnd OAI21X1_526/C vdd NAND2X1
XNAND2X1_499 BUFX4_48/Y operand_A[56] gnd OAI21X1_576/C vdd NAND2X1
XNAND2X1_422 BUFX4_73/Y INVX1_188/Y gnd OAI21X1_457/C vdd NAND2X1
XNAND2X1_455 MUX2X1_62/S OAI21X1_558/B gnd OAI21X1_513/C vdd NAND2X1
XNAND2X1_477 NOR2X1_80/A OAI21X1_333/Y gnd NAND2X1_477/Y vdd NAND2X1
XOAI21X1_950 AOI22X1_58/Y NOR2X1_509/Y NOR2X1_510/Y gnd OAI21X1_950/Y vdd OAI21X1
XINVX2_80 operand_A[55] gnd INVX2_80/Y vdd INVX2
XINVX2_91 INVX2_91/A gnd INVX2_91/Y vdd INVX2
XFILL_31_4_0 gnd vdd FILL
XOAI21X1_21 operand_B[27] operand_A[27] OAI21X1_21/C gnd OAI21X1_22/C vdd OAI21X1
XOAI21X1_76 BUFX4_71/Y OAI21X1_76/B OAI21X1_76/C gnd OAI21X1_76/Y vdd OAI21X1
XOAI21X1_43 INVX2_32/Y MUX2X1_3/S OAI21X1_43/C gnd INVX1_39/A vdd OAI21X1
XOAI21X1_65 XOR2X1_3/A INVX1_47/Y OAI21X1_65/C gnd OAI21X1_66/B vdd OAI21X1
XOAI21X1_87 MUX2X1_23/S XOR2X1_7/A operand_A[63] gnd OAI21X1_88/C vdd OAI21X1
XOAI21X1_54 BUFX4_76/Y OAI21X1_54/B OAI21X1_54/C gnd MUX2X1_2/A vdd OAI21X1
XOAI21X1_32 OAI21X1_32/A OAI21X1_32/B OAI21X1_32/C gnd OAI21X1_32/Y vdd OAI21X1
XOAI21X1_10 INVX1_81/A NOR2X1_21/Y OAI21X1_10/C gnd NOR2X1_24/A vdd OAI21X1
XOAI21X1_98 INVX4_4/Y MUX2X1_3/S OAI21X1_98/C gnd INVX1_60/A vdd OAI21X1
XFILL_22_4_0 gnd vdd FILL
XAND2X2_13 AND2X2_13/A NAND3X1_9/Y gnd AND2X2_13/Y vdd AND2X2
XOAI21X1_257 INVX2_60/Y BUFX4_43/Y OAI21X1_77/C gnd OAI21X1_257/Y vdd OAI21X1
XOAI21X1_202 OAI22X1_3/C NOR2X1_103/A AOI22X1_4/Y gnd OR2X2_4/A vdd OAI21X1
XOAI21X1_224 BUFX4_71/Y MUX2X1_18/Y OAI21X1_224/C gnd INVX1_134/A vdd OAI21X1
XOAI21X1_246 BUFX4_131/Y OAI21X1_76/Y OAI21X1_246/C gnd MUX2X1_120/B vdd OAI21X1
XOAI21X1_268 MUX2X1_87/S OAI21X1_272/A OAI21X1_268/C gnd OAI21X1_268/Y vdd OAI21X1
XOAI21X1_235 INVX4_10/Y BUFX4_67/Y OAI21X1_312/A gnd INVX1_107/A vdd OAI21X1
XOAI21X1_279 INVX1_122/Y MUX2X1_2/S OAI21X1_279/C gnd INVX1_123/A vdd OAI21X1
XOAI21X1_213 XOR2X1_4/A OAI21X1_213/B OAI21X1_213/C gnd OAI21X1_213/Y vdd OAI21X1
XAND2X2_35 operand_A[55] operand_B[55] gnd AND2X2_35/Y vdd AND2X2
XAND2X2_24 OR2X2_24/A OR2X2_24/B gnd AND2X2_24/Y vdd AND2X2
XNAND2X1_252 NOR2X1_54/A MUX2X1_15/Y gnd OAI21X1_223/C vdd NAND2X1
XNAND2X1_230 BUFX4_70/Y INVX1_41/A gnd OAI21X1_197/C vdd NAND2X1
XAND2X2_46 AND2X2_46/A AND2X2_46/B gnd AND2X2_46/Y vdd AND2X2
XNAND2X1_241 BUFX4_74/Y OAI21X1_113/Y gnd OAI21X1_210/C vdd NAND2X1
XAND2X2_57 AND2X2_57/A BUFX4_113/Y gnd AND2X2_57/Y vdd AND2X2
XAND2X2_68 AND2X2_68/A BUFX4_100/Y gnd AND2X2_68/Y vdd AND2X2
XNAND2X1_274 BUFX4_16/Y OAI21X1_405/B gnd OAI21X1_251/C vdd NAND2X1
XNAND2X1_263 BUFX4_69/Y OAI21X1_125/B gnd OAI21X1_312/A vdd NAND2X1
XNAND2X1_296 OR2X2_43/B INVX1_119/Y gnd OAI21X1_273/C vdd NAND2X1
XFILL_5_5_0 gnd vdd FILL
XNAND2X1_285 OR2X2_39/B NOR2X1_141/Y gnd INVX1_209/A vdd NAND2X1
XFILL_13_4_0 gnd vdd FILL
XOAI21X1_791 OAI21X1_791/A OAI21X1_791/B BUFX4_97/Y gnd OAI21X1_792/C vdd OAI21X1
XOAI21X1_780 OAI21X1_780/A BUFX4_77/Y OAI21X1_780/C gnd OAI21X1_780/Y vdd OAI21X1
XINVX1_118 INVX1_118/A gnd INVX1_118/Y vdd INVX1
XINVX1_107 INVX1_107/A gnd INVX1_107/Y vdd INVX1
XINVX1_129 INVX1_129/A gnd INVX1_129/Y vdd INVX1
XNOR2X1_509 NOR2X1_509/A NOR2X1_509/B gnd NOR2X1_509/Y vdd NOR2X1
XINVX4_15 INVX4_15/A gnd INVX4_15/Y vdd INVX4
XINVX4_26 INVX4_26/A gnd INVX4_26/Y vdd INVX4
XFILL_27_3_0 gnd vdd FILL
XFILL_2_3_0 gnd vdd FILL
XFILL_10_2_0 gnd vdd FILL
XNOR2X1_306 NOR2X1_306/A NOR2X1_321/A gnd INVX2_81/A vdd NOR2X1
XFILL_18_3_0 gnd vdd FILL
XNOR2X1_328 INVX4_9/Y INVX2_83/Y gnd INVX1_241/A vdd NOR2X1
XNOR2X1_339 INVX1_244/A INVX1_243/A gnd OR2X2_34/B vdd NOR2X1
XNOR2X1_317 BUFX4_183/Y NOR2X1_317/B gnd INVX1_234/A vdd NOR2X1
XNAND3X1_35 BUFX4_143/Y NAND3X1_35/B NAND3X1_35/C gnd NAND3X1_35/Y vdd NAND3X1
XNOR2X1_46 INVX4_1/A INVX1_26/A gnd NOR2X1_94/B vdd NOR2X1
XNAND3X1_13 INVX1_145/Y OR2X2_14/Y NOR2X1_171/Y gnd NAND3X1_13/Y vdd NAND3X1
XNAND3X1_24 NAND3X1_24/A NAND3X1_24/B NAND3X1_24/C gnd NAND3X1_24/Y vdd NAND3X1
XNOR2X1_24 NOR2X1_24/A NOR2X1_24/B gnd NOR2X1_24/Y vdd NOR2X1
XNOR2X1_35 INVX2_23/Y INVX2_22/Y gnd NOR2X1_35/Y vdd NOR2X1
XNAND3X1_57 BUFX4_97/Y NAND3X1_57/B NAND3X1_57/C gnd NAND3X1_57/Y vdd NAND3X1
XNAND3X1_46 INVX1_266/Y INVX1_267/Y NOR2X1_398/Y gnd NOR2X1_400/A vdd NAND3X1
XNAND3X1_68 NAND3X1_68/A AND2X2_65/Y NAND3X1_68/C gnd NAND3X1_68/Y vdd NAND3X1
XNOR2X1_13 operand_B[17] INVX4_6/Y gnd OAI21X1_7/B vdd NOR2X1
XNOR2X1_68 operand_B[25] INVX4_8/Y gnd NOR2X1_68/Y vdd NOR2X1
XNOR2X1_79 INVX2_36/Y INVX1_51/Y gnd BUFX4_91/A vdd NOR2X1
XNOR2X1_57 OR2X2_7/B INVX4_7/Y gnd NOR2X1_57/Y vdd NOR2X1
XNOR2X1_136 BUFX4_28/Y AND2X2_12/Y gnd NOR2X1_136/Y vdd NOR2X1
XNOR2X1_158 NOR2X1_158/A INVX1_283/A gnd INVX1_127/A vdd NOR2X1
XNOR2X1_103 NOR2X1_103/A INVX4_15/Y gnd AOI22X1_4/C vdd NOR2X1
XMUX2X1_53 MUX2X1_56/B MUX2X1_53/B BUFX4_75/Y gnd MUX2X1_60/B vdd MUX2X1
XMUX2X1_20 MUX2X1_20/A MUX2X1_20/B MUX2X1_71/S gnd MUX2X1_20/Y vdd MUX2X1
XNOR2X1_114 XOR2X1_5/Y OAI21X1_10/C gnd NOR2X1_114/Y vdd NOR2X1
XMUX2X1_86 MUX2X1_97/A MUX2X1_98/B BUFX4_66/Y gnd MUX2X1_87/A vdd MUX2X1
XMUX2X1_97 MUX2X1_97/A MUX2X1_97/B MUX2X1_97/S gnd MUX2X1_99/B vdd MUX2X1
XNOR2X1_147 BUFX4_136/Y NOR2X1_147/B gnd NOR2X1_147/Y vdd NOR2X1
XMUX2X1_31 MUX2X1_31/A MUX2X1_31/B BUFX4_20/Y gnd MUX2X1_32/B vdd MUX2X1
XMUX2X1_75 MUX2X1_75/A MUX2X1_75/B BUFX4_24/Y gnd MUX2X1_75/Y vdd MUX2X1
XMUX2X1_64 MUX2X1_64/A MUX2X1_64/B MUX2X1_64/S gnd MUX2X1_64/Y vdd MUX2X1
XNOR2X1_125 INVX8_4/A INVX8_7/Y gnd BUFX4_87/A vdd NOR2X1
XMUX2X1_42 MUX2X1_42/A MUX2X1_42/B MUX2X1_49/S gnd MUX2X1_42/Y vdd MUX2X1
XNOR2X1_169 operand_B[37] INVX2_55/Y gnd NOR2X1_169/Y vdd NOR2X1
XOAI21X1_609 OAI21X1_623/A INVX2_88/A NOR2X1_359/Y gnd OAI21X1_609/Y vdd OAI21X1
XDFFSR_1 DFFSR_1/Q DFFSR_1/CLK DFFSR_1/R vdd DFFSR_1/D gnd vdd DFFSR
XMUX2X1_109 NOR2X1_470/B MUX2X1_109/B BUFX4_36/Y gnd MUX2X1_109/Y vdd MUX2X1
XNAND2X1_648 operand_B[27] operand_A[27] gnd OAI21X1_935/B vdd NAND2X1
XINVX1_49 INVX1_49/A gnd INVX1_49/Y vdd INVX1
XINVX1_27 INVX1_27/A gnd INVX1_27/Y vdd INVX1
XNAND2X1_637 BUFX4_112/Y OAI21X1_538/C gnd OAI22X1_31/D vdd NAND2X1
XINVX1_16 operand_B[14] gnd INVX1_16/Y vdd INVX1
XNAND2X1_604 AOI22X1_36/Y OAI21X1_782/Y gnd OAI21X1_791/B vdd NAND2X1
XNAND2X1_626 NAND2X1_626/A AOI22X1_44/Y gnd NAND2X1_626/Y vdd NAND2X1
XINVX1_290 INVX1_290/A gnd INVX1_290/Y vdd INVX1
XINVX1_38 INVX1_38/A gnd INVX1_38/Y vdd INVX1
XNAND2X1_615 BUFX4_24/Y OR2X2_39/A gnd OAI21X1_826/C vdd NAND2X1
XFILL_24_1_0 gnd vdd FILL
XNAND2X1_90 BUFX4_67/Y INVX1_93/A gnd OAI21X1_41/C vdd NAND2X1
XAOI21X1_250 NOR2X1_341/A INVX2_86/Y NOR2X1_349/Y gnd OAI21X1_601/C vdd AOI21X1
XAOI21X1_272 NAND3X1_37/Y AOI21X1_272/B NOR2X1_369/Y gnd DFFPOSX1_63/D vdd AOI21X1
XAOI21X1_294 operand_B[63] INVX4_10/Y alu_op[1] gnd AND2X2_50/B vdd AOI21X1
XAOI21X1_261 BUFX4_80/Y NOR2X1_509/A OAI21X1_618/Y gnd NAND3X1_36/B vdd AOI21X1
XAOI21X1_283 INVX1_4/A OAI21X1_650/Y NOR2X1_48/A gnd OAI21X1_651/A vdd AOI21X1
XFILL_7_2_0 gnd vdd FILL
XFILL_15_1_0 gnd vdd FILL
XOAI21X1_428 OR2X2_44/A OR2X2_44/B INVX4_20/A gnd NAND3X1_22/A vdd OAI21X1
XOAI21X1_406 AOI21X1_71/Y BUFX4_35/Y INVX2_48/Y gnd OAI21X1_406/Y vdd OAI21X1
XOAI21X1_417 NOR2X1_147/B BUFX4_136/Y BUFX4_37/Y gnd OAI21X1_418/C vdd OAI21X1
XOAI21X1_439 BUFX4_35/Y INVX1_139/A OAI21X1_439/C gnd MUX2X1_64/A vdd OAI21X1
XNAND2X1_434 OAI21X1_424/Y NOR2X1_244/Y gnd NAND3X1_29/C vdd NAND2X1
XNAND2X1_445 MUX2X1_97/S OAI21X1_467/Y gnd OAI21X1_492/C vdd NAND2X1
XNAND2X1_401 BUFX4_39/Y OAI21X1_301/Y gnd OAI21X1_426/C vdd NAND2X1
XNAND2X1_423 BUFX4_19/Y MUX2X1_52/A gnd OAI21X1_458/C vdd NAND2X1
XNAND2X1_412 NOR2X1_75/A MUX2X1_64/A gnd NAND2X1_417/A vdd NAND2X1
XNAND2X1_489 NOR2X1_310/Y NOR2X1_292/Y gnd NOR2X1_312/A vdd NAND2X1
XNAND2X1_467 MUX2X1_66/S OAI21X1_526/Y gnd OAI21X1_527/C vdd NAND2X1
XNAND2X1_456 BUFX4_18/Y MUX2X1_58/B gnd OAI21X1_514/C vdd NAND2X1
XNAND2X1_478 BUFX4_184/Y OAI21X1_339/Y gnd OAI21X1_548/C vdd NAND2X1
XOAI21X1_940 operand_B[28] operand_A[28] BUFX4_6/Y gnd OAI21X1_941/C vdd OAI21X1
XINVX2_70 operand_B[39] gnd INVX2_70/Y vdd INVX2
XINVX2_81 INVX2_81/A gnd INVX2_81/Y vdd INVX2
XINVX2_92 INVX2_92/A gnd INVX2_92/Y vdd INVX2
XOAI21X1_11 NOR2X1_22/Y NOR2X1_23/Y NAND3X1_4/B gnd NOR2X1_24/B vdd OAI21X1
XFILL_31_4_1 gnd vdd FILL
XOAI21X1_77 INVX2_45/Y MUX2X1_3/S OAI21X1_77/C gnd OAI21X1_77/Y vdd OAI21X1
XOAI21X1_33 operand_B[27] INVX2_30/Y OAI21X1_33/C gnd AOI22X1_1/B vdd OAI21X1
XOAI21X1_22 OR2X2_2/A OAI21X1_22/B OAI21X1_22/C gnd INVX1_25/A vdd OAI21X1
XOAI21X1_44 INVX2_31/Y BUFX4_43/Y OAI21X1_44/C gnd INVX1_95/A vdd OAI21X1
XOAI21X1_88 INVX1_52/Y INVX8_3/A OAI21X1_88/C gnd INVX1_53/A vdd OAI21X1
XOAI21X1_66 BUFX4_134/Y OAI21X1_66/B OAI21X1_66/C gnd OR2X2_13/A vdd OAI21X1
XOAI21X1_55 INVX2_21/Y BUFX4_43/Y OAI21X1_55/C gnd OAI21X1_55/Y vdd OAI21X1
XOAI21X1_99 INVX2_8/Y BUFX4_43/Y OAI21X1_99/C gnd OAI21X1_99/Y vdd OAI21X1
XFILL_22_4_1 gnd vdd FILL
XOAI21X1_203 MUX2X1_25/Y INVX8_15/Y AOI21X1_63/Y gnd OR2X2_5/B vdd OAI21X1
XAND2X2_36 AND2X2_36/A AND2X2_36/B gnd AND2X2_36/Y vdd AND2X2
XOAI21X1_258 INVX1_97/Y BUFX4_75/Y OAI21X1_258/C gnd INVX1_115/A vdd OAI21X1
XAND2X2_14 AND2X2_14/A BUFX4_159/Y gnd AND2X2_14/Y vdd AND2X2
XOAI21X1_247 OAI21X1_247/A BUFX4_21/Y OAI21X1_247/C gnd MUX2X1_124/B vdd OAI21X1
XOAI21X1_225 BUFX4_122/Y OAI21X1_225/B OAI21X1_225/C gnd OAI21X1_228/A vdd OAI21X1
XOAI21X1_269 BUFX4_39/Y MUX2X1_39/B OAI21X1_269/C gnd AOI21X1_78/B vdd OAI21X1
XOAI21X1_236 INVX1_107/Y BUFX4_120/Y OAI21X1_236/C gnd MUX2X1_29/A vdd OAI21X1
XAND2X2_25 AND2X2_25/A BUFX4_184/Y gnd OAI22X1_8/C vdd AND2X2
XAND2X2_47 AND2X2_47/A NOR2X1_56/Y gnd AND2X2_47/Y vdd AND2X2
XOAI21X1_214 INVX1_61/Y BUFX4_192/Y OAI21X1_214/C gnd INVX1_104/A vdd OAI21X1
XNAND2X1_231 operand_A[31] BUFX4_53/Y gnd OAI21X1_198/C vdd NAND2X1
XNAND2X1_253 BUFX4_71/Y OAI21X1_135/Y gnd OAI21X1_224/C vdd NAND2X1
XNAND2X1_275 BUFX4_134/Y INVX1_52/A gnd OAI21X1_249/C vdd NAND2X1
XNAND2X1_286 INVX4_18/A NOR2X1_142/Y gnd NAND3X1_10/C vdd NAND2X1
XNAND2X1_264 NOR2X1_75/A OAI21X1_234/Y gnd AOI21X1_66/B vdd NAND2X1
XNAND2X1_220 NOR2X1_54/A MUX2X1_4/Y gnd OAI21X1_187/C vdd NAND2X1
XNAND2X1_242 NOR2X1_54/A MUX2X1_11/Y gnd OAI21X1_211/C vdd NAND2X1
XFILL_5_5_1 gnd vdd FILL
XAND2X2_58 AND2X2_58/A AND2X2_58/B gnd AND2X2_58/Y vdd AND2X2
XAND2X2_69 OR2X2_7/A MUX2X1_34/S gnd AND2X2_69/Y vdd AND2X2
XFILL_29_0_0 gnd vdd FILL
XFILL_4_0_0 gnd vdd FILL
XNAND2X1_297 INVX8_3/A OAI21X1_100/Y gnd OAI21X1_274/C vdd NAND2X1
XFILL_13_4_1 gnd vdd FILL
XOAI21X1_781 OAI21X1_781/A XNOR2X1_19/Y INVX1_303/Y gnd OAI21X1_782/B vdd OAI21X1
XOAI21X1_792 BUFX4_97/Y INVX1_304/Y OAI21X1_792/C gnd DFFPOSX1_8/D vdd OAI21X1
XOAI21X1_770 BUFX4_184/Y OAI21X1_770/B NOR2X1_447/Y gnd OAI21X1_780/C vdd OAI21X1
XINVX1_108 INVX1_108/A gnd INVX1_108/Y vdd INVX1
XINVX1_119 INVX1_119/A gnd INVX1_119/Y vdd INVX1
XFILL_4_1 gnd vdd FILL
XINVX4_16 INVX4_16/A gnd INVX4_16/Y vdd INVX4
XFILL_27_3_1 gnd vdd FILL
XFILL_2_3_1 gnd vdd FILL
XFILL_10_2_1 gnd vdd FILL
XNOR2X1_307 NOR2X1_307/A NOR2X1_307/B gnd NOR2X1_307/Y vdd NOR2X1
XNOR2X1_329 NOR2X1_333/A INVX1_241/A gnd INVX2_84/A vdd NOR2X1
XNOR2X1_318 INVX4_13/Y INVX1_235/Y gnd NOR2X1_320/B vdd NOR2X1
XFILL_18_3_1 gnd vdd FILL
XAOI21X1_410 OAI21X1_937/Y NOR2X1_506/Y NOR2X1_507/Y gnd DFFPOSX1_29/D vdd AOI21X1
XNAND3X1_14 MUX2X1_64/S OR2X2_39/B INVX1_66/A gnd NAND3X1_14/Y vdd NAND3X1
XNOR2X1_47 BUFX4_29/Y NOR2X1_94/B gnd NOR2X1_47/Y vdd NOR2X1
XNOR2X1_69 operand_B[24] INVX2_32/Y gnd NOR2X1_69/Y vdd NOR2X1
XNAND3X1_36 NAND3X1_36/A NAND3X1_36/B NAND3X1_36/C gnd NAND3X1_36/Y vdd NAND3X1
XNAND3X1_25 NAND3X1_25/A OR2X2_25/Y NAND3X1_25/C gnd NAND3X1_25/Y vdd NAND3X1
XNAND3X1_69 NAND3X1_69/A NAND3X1_69/B NAND3X1_69/C gnd NOR2X1_479/B vdd NAND3X1
XNAND3X1_47 INVX1_268/Y INVX1_269/Y NOR2X1_399/Y gnd NOR2X1_400/B vdd NAND3X1
XNOR2X1_36 INVX2_20/Y INVX1_18/Y gnd NOR2X1_36/Y vdd NOR2X1
XNOR2X1_25 INVX1_13/Y INVX1_12/Y gnd NOR2X1_25/Y vdd NOR2X1
XNOR2X1_58 operand_B[6] INVX2_13/Y gnd NOR2X1_58/Y vdd NOR2X1
XNAND3X1_58 NAND3X1_58/A NAND3X1_58/B NAND3X1_58/C gnd NOR2X1_433/A vdd NAND3X1
XNOR2X1_14 OAI21X1_3/A OAI21X1_7/Y gnd AND2X2_1/B vdd NOR2X1
XNOR2X1_137 operand_B[32] INVX2_45/Y gnd NOR2X1_137/Y vdd NOR2X1
XNOR2X1_104 OR2X2_2/A OR2X2_2/B gnd NOR2X1_104/Y vdd NOR2X1
XMUX2X1_10 operand_A[63] operand_A[62] BUFX4_48/Y gnd NOR2X1_82/B vdd MUX2X1
XMUX2X1_65 MUX2X1_65/A MUX2X1_65/B BUFX4_75/Y gnd MUX2X1_66/A vdd MUX2X1
XNOR2X1_148 OR2X2_8/B NOR2X1_148/B gnd NOR2X1_148/Y vdd NOR2X1
XMUX2X1_54 MUX2X1_54/A MUX2X1_54/B BUFX4_39/Y gnd MUX2X1_54/Y vdd MUX2X1
XMUX2X1_21 MUX2X1_21/A MUX2X1_21/B OR2X2_43/B gnd MUX2X1_21/Y vdd MUX2X1
XMUX2X1_43 MUX2X1_55/A MUX2X1_43/B BUFX4_25/Y gnd MUX2X1_44/A vdd MUX2X1
XNOR2X1_115 NAND3X1_1/A OR2X2_45/B gnd NOR2X1_115/Y vdd NOR2X1
XNOR2X1_126 NOR2X1_82/A INVX2_58/Y gnd INVX1_98/A vdd NOR2X1
XMUX2X1_76 MUX2X1_76/A MUX2X1_76/B BUFX4_74/Y gnd MUX2X1_76/Y vdd MUX2X1
XMUX2X1_98 MUX2X1_98/A MUX2X1_98/B MUX2X1_98/S gnd MUX2X1_99/A vdd MUX2X1
XMUX2X1_87 MUX2X1_87/A MUX2X1_87/B MUX2X1_87/S gnd MUX2X1_95/B vdd MUX2X1
XNOR2X1_159 BUFX4_42/Y OR2X2_22/A gnd INVX1_132/A vdd NOR2X1
XMUX2X1_32 MUX2X1_32/A MUX2X1_32/B MUX2X1_32/S gnd OAI22X1_4/C vdd MUX2X1
XNAND2X1_605 MUX2X1_99/S OAI21X1_734/B gnd OAI21X1_784/C vdd NAND2X1
XINVX1_280 INVX1_280/A gnd INVX1_280/Y vdd INVX1
XINVX1_291 INVX1_291/A gnd INVX1_291/Y vdd INVX1
XNAND2X1_616 BUFX4_36/Y OAI21X1_738/B gnd OAI21X1_827/C vdd NAND2X1
XNAND2X1_627 OR2X2_46/B BUFX4_152/Y gnd AND2X2_66/B vdd NAND2X1
XNAND2X1_649 NOR2X1_503/Y OAI22X1_37/Y gnd NAND2X1_649/Y vdd NAND2X1
XINVX1_28 INVX1_28/A gnd INVX1_28/Y vdd INVX1
XNAND2X1_638 NOR2X1_495/Y OAI22X1_31/Y gnd NAND2X1_638/Y vdd NAND2X1
XINVX1_17 INVX1_17/A gnd INVX1_17/Y vdd INVX1
XNAND2X1_91 BUFX4_119/Y INVX1_113/A gnd OAI21X1_42/C vdd NAND2X1
XNAND2X1_80 INVX4_26/A XNOR2X1_25/Y gnd NOR2X1_66/B vdd NAND2X1
XINVX1_39 INVX1_39/A gnd INVX1_39/Y vdd INVX1
XFILL_24_1_1 gnd vdd FILL
XAOI21X1_240 OR2X2_34/B OR2X2_34/A BUFX4_30/Y gnd AOI21X1_245/A vdd AOI21X1
XAOI21X1_251 INVX1_248/Y OAI21X1_566/B INVX1_253/A gnd OAI21X1_623/A vdd AOI21X1
XAOI21X1_273 INVX4_25/Y OAI21X1_627/Y BUFX4_94/Y gnd AOI21X1_275/B vdd AOI21X1
XAOI21X1_262 AOI21X1_262/A OAI21X1_609/Y NAND3X1_36/Y gnd AOI21X1_263/A vdd AOI21X1
XAOI21X1_284 operand_B[29] INVX2_2/Y NOR2X1_414/Y gnd OAI21X1_654/A vdd AOI21X1
XAOI21X1_295 OAI21X1_655/Y NOR2X1_424/Y alu_op[0] gnd OAI21X1_675/A vdd AOI21X1
XFILL_7_2_1 gnd vdd FILL
XFILL_15_1_1 gnd vdd FILL
XOAI21X1_407 OAI22X1_7/C NOR2X1_202/A AOI22X1_11/Y gnd OR2X2_20/A vdd OAI21X1
XOAI21X1_418 INVX1_123/A BUFX4_38/Y OAI21X1_418/C gnd OAI22X1_19/A vdd OAI21X1
XOAI21X1_429 INVX8_2/A MUX2X1_31/B OR2X2_22/Y gnd INVX1_177/A vdd OAI21X1
XNAND2X1_435 NOR2X1_245/Y INVX1_198/Y gnd OAI21X1_472/B vdd NAND2X1
XNAND2X1_413 BUFX4_46/Y operand_A[44] gnd OAI21X1_440/C vdd NAND2X1
XNAND2X1_446 MUX2X1_99/S OAI21X1_441/Y gnd OAI21X1_493/C vdd NAND2X1
XNAND2X1_402 INVX4_18/A INVX1_310/A gnd NAND3X1_22/C vdd NAND2X1
XNAND2X1_457 INVX2_49/A AOI21X1_78/B gnd OAI21X1_515/C vdd NAND2X1
XNAND2X1_468 MUX2X1_34/S MUX2X1_32/A gnd OAI21X1_528/C vdd NAND2X1
XNAND2X1_424 MUX2X1_32/S INVX1_261/A gnd OAI21X1_459/C vdd NAND2X1
XNAND2X1_479 BUFX4_186/Y NOR2X1_170/B gnd OAI21X1_549/C vdd NAND2X1
XOAI21X1_941 BUFX4_63/Y INVX1_327/Y OAI21X1_941/C gnd NOR2X1_505/B vdd OAI21X1
XOAI21X1_930 INVX1_325/Y XNOR2X1_27/Y OAI21X1_20/C gnd OAI21X1_931/B vdd OAI21X1
XNOR2X1_490 NOR2X1_490/A NOR2X1_490/B gnd NOR2X1_490/Y vdd NOR2X1
XINVX2_82 INVX2_82/A gnd INVX2_82/Y vdd INVX2
XINVX2_60 operand_A[34] gnd INVX2_60/Y vdd INVX2
XINVX2_71 operand_A[42] gnd INVX2_71/Y vdd INVX2
XINVX2_93 INVX2_93/A gnd INVX2_93/Y vdd INVX2
XOAI21X1_23 OAI21X1_23/A OR2X2_2/Y INVX1_25/Y gnd AND2X2_74/A vdd OAI21X1
XOAI21X1_34 OAI21X1_34/A INVX1_33/Y AOI22X1_1/Y gnd OAI21X1_34/Y vdd OAI21X1
XOAI21X1_12 BUFX4_82/Y INVX2_14/Y OAI21X1_12/C gnd OAI21X1_13/C vdd OAI21X1
XOAI21X1_45 INVX1_39/Y BUFX4_67/Y OAI21X1_45/C gnd INVX1_40/A vdd OAI21X1
XOAI21X1_67 INVX2_40/Y MUX2X1_8/S OAI21X1_67/C gnd OAI21X1_69/B vdd OAI21X1
XOAI21X1_78 BUFX4_190/Y MUX2X1_7/Y OAI21X1_78/C gnd INVX1_293/A vdd OAI21X1
XOAI21X1_89 INVX1_53/Y BUFX4_42/Y INVX2_48/Y gnd INVX1_54/A vdd OAI21X1
XOAI21X1_56 BUFX4_192/Y MUX2X1_3/Y OAI21X1_56/C gnd INVX1_45/A vdd OAI21X1
XOAI21X1_204 INVX1_78/Y INVX4_15/Y INVX4_16/Y gnd NAND3X1_6/C vdd OAI21X1
XOAI21X1_226 BUFX4_71/Y MUX2X1_17/Y OAI21X1_226/C gnd MUX2X1_27/B vdd OAI21X1
XOAI21X1_237 MUX2X1_29/Y BUFX4_164/Y OR2X2_7/Y gnd AND2X2_52/A vdd OAI21X1
XOAI21X1_215 INVX1_60/Y MUX2X1_98/S OAI21X1_215/C gnd OAI21X1_215/Y vdd OAI21X1
XAND2X2_26 AND2X2_26/A AND2X2_26/B gnd AND2X2_26/Y vdd AND2X2
XAND2X2_15 AND2X2_15/A AND2X2_15/B gnd AND2X2_15/Y vdd AND2X2
XAND2X2_37 AND2X2_37/A AND2X2_37/B gnd AND2X2_37/Y vdd AND2X2
XOAI21X1_248 BUFX4_133/Y OAI21X1_73/A OAI21X1_248/C gnd OAI21X1_405/B vdd OAI21X1
XOAI21X1_259 INVX1_115/Y INVX8_3/A OAI21X1_259/C gnd MUX2X1_38/A vdd OAI21X1
XAND2X2_48 AND2X2_48/A AND2X2_48/B gnd AND2X2_48/Y vdd AND2X2
XAND2X2_59 AND2X2_59/A BUFX4_116/Y gnd AND2X2_59/Y vdd AND2X2
XFILL_29_0_1 gnd vdd FILL
XNAND2X1_287 INVX2_61/Y INVX1_116/Y gnd AOI22X1_6/D vdd NAND2X1
XNAND2X1_232 MUX2X1_97/S OAI21X1_47/Y gnd OAI21X1_199/C vdd NAND2X1
XNAND2X1_298 BUFX4_68/Y OAI21X1_275/Y gnd OAI21X1_276/C vdd NAND2X1
XNAND2X1_210 MUX2X1_30/S OAI21X1_176/Y gnd OAI21X1_177/C vdd NAND2X1
XNAND2X1_254 MUX2X1_71/S INVX1_134/A gnd OAI21X1_225/C vdd NAND2X1
XNAND2X1_265 BUFX4_83/Y AOI21X1_66/Y gnd NAND3X1_8/A vdd NAND2X1
XNAND2X1_276 BUFX4_183/Y OAI21X1_250/Y gnd AOI21X1_72/B vdd NAND2X1
XNAND2X1_243 NOR2X1_19/B MUX2X1_35/B gnd OAI21X1_212/C vdd NAND2X1
XNAND2X1_221 MUX2X1_99/S OAI21X1_187/Y gnd OAI21X1_189/C vdd NAND2X1
XFILL_4_0_1 gnd vdd FILL
XOAI21X1_782 XOR2X1_5/Y OAI21X1_782/B OAI21X1_782/C gnd OAI21X1_782/Y vdd OAI21X1
XOAI21X1_793 AOI21X1_9/Y INVX1_17/A BUFX4_105/Y gnd OAI21X1_793/Y vdd OAI21X1
XOAI21X1_760 XOR2X1_7/A MUX2X1_94/B OAI21X1_760/C gnd NOR2X1_470/B vdd OAI21X1
XOAI21X1_771 OR2X2_14/A BUFX4_77/Y OAI21X1_780/C gnd OAI21X1_771/Y vdd OAI21X1
XINVX1_109 INVX1_109/A gnd INVX1_109/Y vdd INVX1
XOAI21X1_590 INVX4_9/Y INVX2_83/Y OAI21X1_590/C gnd OR2X2_34/A vdd OAI21X1
XFILL_4_2 gnd vdd FILL
XINVX4_17 INVX4_17/A gnd INVX4_17/Y vdd INVX4
XNOR2X1_308 INVX2_81/Y INVX1_232/A gnd NOR2X1_321/B vdd NOR2X1
XNOR2X1_319 operand_A[57] operand_B[57] gnd NOR2X1_320/A vdd NOR2X1
XAOI21X1_400 BUFX4_81/Y MUX2X1_127/Y INVX8_9/Y gnd OAI22X1_35/C vdd AOI21X1
XAOI21X1_411 NOR2X1_3/A NOR2X1_508/Y BUFX4_29/Y gnd OAI21X1_943/C vdd AOI21X1
XFILL_20_5_0 gnd vdd FILL
XNAND3X1_37 BUFX4_107/Y NAND3X1_38/C NAND3X1_37/C gnd NAND3X1_37/Y vdd NAND3X1
XNAND3X1_26 INVX4_22/Y INVX1_192/Y NAND3X1_26/C gnd NAND3X1_27/B vdd NAND3X1
XNAND3X1_15 OR2X2_15/Y NAND3X1_15/B OR2X2_16/Y gnd NAND3X1_15/Y vdd NAND3X1
XNAND3X1_48 INVX1_270/Y INVX1_271/Y NOR2X1_401/Y gnd NOR2X1_403/A vdd NAND3X1
XNOR2X1_48 NOR2X1_48/A NOR2X1_48/B gnd NOR2X1_48/Y vdd NOR2X1
XNOR2X1_37 INVX2_21/Y INVX1_19/Y gnd NOR2X1_37/Y vdd NOR2X1
XNOR2X1_15 BUFX4_66/Y INVX2_9/Y gnd NOR2X1_15/Y vdd NOR2X1
XNOR2X1_59 NOR2X1_59/A INVX1_82/A gnd NOR2X1_59/Y vdd NOR2X1
XNOR2X1_26 INVX2_13/Y INVX1_14/Y gnd NOR2X1_26/Y vdd NOR2X1
XNAND3X1_59 NAND3X1_59/A NAND3X1_59/B NOR2X1_437/Y gnd NOR2X1_438/B vdd NAND3X1
XFILL_11_5_0 gnd vdd FILL
XMUX2X1_11 operand_A[6] operand_A[7] MUX2X1_8/S gnd MUX2X1_11/Y vdd MUX2X1
XNOR2X1_105 INVX4_1/A OAI21X1_94/C gnd AND2X2_9/A vdd NOR2X1
XNOR2X1_138 operand_B[33] INVX2_56/Y gnd NOR2X1_138/Y vdd NOR2X1
XMUX2X1_77 operand_A[30] operand_A[29] MUX2X1_1/S gnd MUX2X1_77/Y vdd MUX2X1
XMUX2X1_22 MUX2X1_22/A MUX2X1_22/B BUFX4_69/Y gnd MUX2X1_22/Y vdd MUX2X1
XMUX2X1_66 MUX2X1_66/A MUX2X1_66/B MUX2X1_66/S gnd MUX2X1_67/B vdd MUX2X1
XMUX2X1_33 MUX2X1_33/A MUX2X1_33/B INVX8_2/A gnd MUX2X1_33/Y vdd MUX2X1
XMUX2X1_55 MUX2X1_55/A MUX2X1_55/B OR2X2_13/B gnd MUX2X1_55/Y vdd MUX2X1
XMUX2X1_44 MUX2X1_44/A MUX2X1_44/B MUX2X1_49/S gnd MUX2X1_44/Y vdd MUX2X1
XNOR2X1_149 NOR2X1_149/A NOR2X1_149/B gnd NOR2X1_149/Y vdd NOR2X1
XNOR2X1_116 XOR2X1_6/Y XOR2X1_8/Y gnd NOR2X1_116/Y vdd NOR2X1
XMUX2X1_88 operand_A[16] operand_A[15] MUX2X1_5/S gnd MUX2X1_90/B vdd MUX2X1
XMUX2X1_99 MUX2X1_99/A MUX2X1_99/B MUX2X1_99/S gnd MUX2X1_99/Y vdd MUX2X1
XNOR2X1_127 MUX2X1_51/S INVX1_98/Y gnd INVX1_99/A vdd NOR2X1
XNAND2X1_639 INVX1_9/Y INVX4_3/Y gnd AOI22X1_52/D vdd NAND2X1
XNAND2X1_628 OR2X2_47/B OR2X2_47/A gnd NAND3X1_70/B vdd NAND2X1
XINVX1_18 operand_B[13] gnd INVX1_18/Y vdd INVX1
XINVX1_281 INVX1_281/A gnd INVX1_281/Y vdd INVX1
XINVX1_29 operand_A[0] gnd INVX1_29/Y vdd INVX1
XINVX1_292 INVX1_292/A gnd INVX1_292/Y vdd INVX1
XNAND2X1_606 BUFX4_90/Y OAI21X1_786/Y gnd NAND2X1_608/A vdd NAND2X1
XINVX1_270 BUFX2_22/A gnd INVX1_270/Y vdd INVX1
XNAND2X1_617 OR2X2_40/B AOI22X1_12/A gnd OAI21X1_829/C vdd NAND2X1
XNAND2X1_81 NOR2X1_48/Y NOR2X1_66/Y gnd INVX1_31/A vdd NAND2X1
XNAND2X1_92 BUFX4_53/Y operand_A[23] gnd OAI21X1_43/C vdd NAND2X1
XNAND2X1_70 BUFX4_37/Y INVX2_11/Y gnd INVX1_280/A vdd NAND2X1
XAOI21X1_230 OAI21X1_573/Y NOR2X1_325/Y OAI21X1_581/Y gnd AOI21X1_231/A vdd AOI21X1
XAOI21X1_252 INVX2_88/A OAI21X1_623/A OAI21X1_602/Y gnd NOR2X1_352/B vdd AOI21X1
XAOI21X1_241 BUFX4_167/Y MUX2X1_58/Y INVX8_7/Y gnd AOI21X1_243/A vdd AOI21X1
XAOI21X1_263 AOI21X1_263/A OAI21X1_608/Y NOR2X1_363/Y gnd DFFPOSX1_62/D vdd AOI21X1
XAOI21X1_285 INVX1_76/Y OAI21X1_94/C NOR2X1_415/Y gnd OAI21X1_654/C vdd AOI21X1
XAOI21X1_274 XOR2X1_3/A INVX1_254/A OAI21X1_628/Y gnd OAI21X1_629/C vdd AOI21X1
XAOI21X1_296 INVX2_34/Y NOR2X1_413/Y NAND2X1_556/Y gnd OAI21X1_675/C vdd AOI21X1
XOAI21X1_408 INVX2_71/Y INVX2_72/Y OAI21X1_408/C gnd OAI21X1_409/B vdd OAI21X1
XFILL_21_1 gnd vdd FILL
XOAI21X1_419 AND2X2_20/Y INVX2_48/A BUFX4_179/Y gnd OAI21X1_419/Y vdd OAI21X1
XNAND2X1_458 NOR2X1_271/B BUFX4_149/Y gnd NAND3X1_30/A vdd NAND2X1
XNAND2X1_469 NAND2X1_469/A NOR2X1_282/Y gnd OAI21X1_529/B vdd NAND2X1
XNAND2X1_436 INVX1_200/A INVX1_158/Y gnd INVX1_199/A vdd NAND2X1
XNAND2X1_425 operand_A[47] operand_B[47] gnd INVX1_194/A vdd NAND2X1
XNAND2X1_414 BUFX4_191/Y OAI21X1_412/Y gnd OAI21X1_441/C vdd NAND2X1
XNAND2X1_447 INVX8_8/A OAI21X1_213/Y gnd OAI21X1_494/C vdd NAND2X1
XNAND2X1_403 BUFX4_19/Y INVX1_129/A gnd OAI21X1_431/C vdd NAND2X1
XFILL_25_4_0 gnd vdd FILL
XFILL_0_4_0 gnd vdd FILL
XNOR2X1_480 OR2X2_48/A BUFX2_18/A gnd NOR2X1_480/Y vdd NOR2X1
XOAI21X1_942 BUFX4_158/Y NOR2X1_3/B BUFX4_99/Y gnd NOR2X1_505/A vdd OAI21X1
XOAI21X1_931 NOR2X1_67/A OAI21X1_931/B OAI21X1_931/C gnd AOI22X1_57/D vdd OAI21X1
XOAI21X1_920 OR2X2_48/A INVX1_322/Y OAI21X1_920/C gnd OAI21X1_920/Y vdd OAI21X1
XNOR2X1_491 XNOR2X1_13/Y BUFX4_155/Y gnd NOR2X1_492/A vdd NOR2X1
XFILL_8_5_0 gnd vdd FILL
XINVX2_83 operand_B[58] gnd INVX2_83/Y vdd INVX2
XINVX2_50 operand_A[31] gnd INVX2_50/Y vdd INVX2
XINVX2_61 operand_A[35] gnd INVX2_61/Y vdd INVX2
XINVX2_72 operand_B[42] gnd INVX2_72/Y vdd INVX2
XINVX2_94 INVX2_94/A gnd INVX2_94/Y vdd INVX2
XOAI21X1_24 INVX4_1/Y INVX1_26/Y NOR2X1_47/Y gnd OAI21X1_24/Y vdd OAI21X1
XOAI21X1_35 NOR2X1_96/B INVX4_1/Y BUFX4_141/Y gnd OAI21X1_35/Y vdd OAI21X1
XOAI21X1_68 INVX2_41/Y MUX2X1_4/S OAI21X1_68/C gnd INVX1_48/A vdd OAI21X1
XOAI21X1_46 INVX4_2/Y MUX2X1_9/S OAI21X1_46/C gnd INVX1_41/A vdd OAI21X1
XFILL_16_4_0 gnd vdd FILL
XOAI21X1_57 INVX2_26/Y BUFX4_46/Y OAI21X1_57/C gnd OAI21X1_57/Y vdd OAI21X1
XOAI21X1_13 BUFX4_111/Y operand_A[5] OAI21X1_13/C gnd OAI21X1_14/B vdd OAI21X1
XOAI21X1_79 BUFX4_136/Y INVX1_293/A OAI21X1_79/C gnd OAI21X1_85/B vdd OAI21X1
XOAI21X1_205 INVX2_45/Y operand_B[32] AOI21X1_64/A gnd XNOR2X1_30/A vdd OAI21X1
XOAI21X1_238 BUFX4_62/Y OAI21X1_239/C AOI22X1_5/Y gnd OR2X2_8/A vdd OAI21X1
XOAI21X1_227 BUFX4_72/Y MUX2X1_19/Y OAI21X1_227/C gnd MUX2X1_27/A vdd OAI21X1
XOAI21X1_249 OAI21X1_62/Y MUX2X1_87/S OAI21X1_249/C gnd INVX1_109/A vdd OAI21X1
XOAI21X1_216 INVX1_104/Y BUFX4_136/Y OAI21X1_216/C gnd MUX2X1_26/B vdd OAI21X1
XAND2X2_49 AND2X2_49/A INVX1_248/Y gnd AND2X2_49/Y vdd AND2X2
XAND2X2_16 INVX1_162/A AND2X2_16/B gnd AND2X2_16/Y vdd AND2X2
XAND2X2_38 AND2X2_38/A AND2X2_38/B gnd AND2X2_38/Y vdd AND2X2
XAND2X2_27 AND2X2_27/A AND2X2_27/B gnd AND2X2_27/Y vdd AND2X2
XNAND2X1_211 INVX8_3/A MUX2X1_23/Y gnd OAI21X1_178/C vdd NAND2X1
XNAND2X1_200 NOR2X1_115/Y INVX1_82/Y gnd OAI21X1_164/A vdd NAND2X1
XNAND2X1_288 operand_A[35] operand_B[35] gnd OAI21X1_283/C vdd NAND2X1
XNAND2X1_255 BUFX4_71/Y OAI21X1_140/Y gnd OAI21X1_226/C vdd NAND2X1
XNAND2X1_233 BUFX4_120/Y OAI21X1_199/Y gnd OAI21X1_200/C vdd NAND2X1
XNAND2X1_266 BUFX4_120/Y MUX2X1_28/B gnd OAI21X1_236/C vdd NAND2X1
XNAND2X1_277 MUX2X1_2/S OAI21X1_58/Y gnd OAI21X1_253/C vdd NAND2X1
XNAND2X1_222 BUFX4_191/Y MUX2X1_3/Y gnd OAI21X1_188/C vdd NAND2X1
XNAND2X1_244 INVX8_2/A INVX1_103/Y gnd OAI21X1_213/C vdd NAND2X1
XNAND2X1_299 MUX2X1_99/S OAI21X1_107/Y gnd OAI21X1_277/C vdd NAND2X1
XOAI21X1_772 AOI21X1_51/Y OR2X2_3/B OAI21X1_29/B gnd INVX1_302/A vdd OAI21X1
XOAI21X1_783 INVX1_302/Y INVX1_281/Y NAND2X1_23/A gnd XNOR2X1_40/A vdd OAI21X1
XOAI21X1_750 NOR2X1_57/Y INVX2_92/Y OAI21X1_9/Y gnd INVX1_297/A vdd OAI21X1
XOAI21X1_794 INVX1_17/A AOI21X1_55/B OAI21X1_794/C gnd OAI21X1_795/C vdd OAI21X1
XOAI21X1_761 MUX2X1_27/S MUX2X1_27/A OAI21X1_761/C gnd INVX1_299/A vdd OAI21X1
XFILL_31_2_0 gnd vdd FILL
XFILL_22_2_0 gnd vdd FILL
XBUFX4_90 BUFX4_91/A gnd BUFX4_90/Y vdd BUFX4
XFILL_5_3_0 gnd vdd FILL
XFILL_13_2_0 gnd vdd FILL
XOAI21X1_591 INVX2_85/Y MUX2X1_6/S OAI21X1_591/C gnd OAI21X1_614/B vdd OAI21X1
XOAI21X1_580 OAI21X1_917/A OR2X2_16/B AND2X2_40/Y gnd OAI21X1_580/Y vdd OAI21X1
XINVX4_18 INVX4_18/A gnd OR2X2_32/B vdd INVX4
XNOR2X1_309 BUFX4_30/Y NOR2X1_321/B gnd NOR2X1_309/Y vdd NOR2X1
XFILL_20_5_1 gnd vdd FILL
XAOI21X1_401 NAND2X1_59/A BUFX4_57/Y NAND2X1_644/Y gnd OAI21X1_918/C vdd AOI21X1
XAOI21X1_412 MUX2X1_64/S INVX1_328/Y BUFX4_111/Y gnd OAI21X1_945/C vdd AOI21X1
XNAND3X1_16 INVX4_19/A INVX2_65/Y NOR2X1_181/Y gnd OR2X2_17/B vdd NAND3X1
XNAND3X1_38 INVX2_91/Y INVX4_25/Y NAND3X1_38/C gnd NAND3X1_39/B vdd NAND3X1
XNAND3X1_27 NAND3X1_9/A NAND3X1_27/B NAND3X1_27/C gnd NAND3X1_27/Y vdd NAND3X1
XNAND3X1_49 INVX1_272/Y INVX1_273/Y NOR2X1_402/Y gnd NOR2X1_403/B vdd NAND3X1
XFILL_27_1_0 gnd vdd FILL
XNOR2X1_27 XNOR2X1_4/Y XNOR2X1_5/Y gnd NOR2X1_27/Y vdd NOR2X1
XFILL_2_1_0 gnd vdd FILL
XNOR2X1_38 operand_A[13] operand_B[13] gnd INVX1_21/A vdd NOR2X1
XNOR2X1_16 OR2X2_39/B INVX2_11/Y gnd NOR2X1_16/Y vdd NOR2X1
XNOR2X1_49 operand_B[16] INVX2_6/Y gnd NOR2X1_49/Y vdd NOR2X1
XFILL_10_0_0 gnd vdd FILL
XFILL_11_5_1 gnd vdd FILL
XNOR2X1_106 NOR2X1_106/A NOR2X1_106/B gnd NOR2X1_106/Y vdd NOR2X1
XMUX2X1_23 NOR2X1_82/B MUX2X1_5/Y MUX2X1_23/S gnd MUX2X1_23/Y vdd MUX2X1
XFILL_18_1_0 gnd vdd FILL
XMUX2X1_45 MUX2X1_51/A MUX2X1_45/B MUX2X1_66/S gnd MUX2X1_45/Y vdd MUX2X1
XMUX2X1_12 operand_A[10] operand_A[11] MUX2X1_9/S gnd MUX2X1_12/Y vdd MUX2X1
XMUX2X1_34 MUX2X1_34/A MUX2X1_34/B MUX2X1_34/S gnd MUX2X1_34/Y vdd MUX2X1
XMUX2X1_56 MUX2X1_59/B MUX2X1_56/B BUFX4_75/Y gnd MUX2X1_66/B vdd MUX2X1
XMUX2X1_78 operand_A[28] operand_A[27] BUFX4_50/Y gnd MUX2X1_78/Y vdd MUX2X1
XNOR2X1_139 INVX4_10/Y BUFX4_69/Y gnd NOR2X1_139/Y vdd NOR2X1
XMUX2X1_67 MUX2X1_67/A MUX2X1_67/B BUFX4_35/Y gnd MUX2X1_67/Y vdd MUX2X1
XNOR2X1_117 operand_A[9] INVX2_25/Y gnd NOR2X1_117/Y vdd NOR2X1
XMUX2X1_89 operand_A[14] operand_A[13] BUFX4_48/Y gnd MUX2X1_90/A vdd MUX2X1
XNOR2X1_128 BUFX4_42/Y INVX1_99/Y gnd NOR2X1_128/Y vdd NOR2X1
XINVX1_260 INVX1_260/A gnd INVX1_260/Y vdd INVX1
XINVX1_293 INVX1_293/A gnd INVX1_293/Y vdd INVX1
XINVX1_19 operand_B[12] gnd INVX1_19/Y vdd INVX1
XNAND2X1_618 NAND2X1_618/A AOI22X1_41/Y gnd NAND2X1_618/Y vdd NAND2X1
XNAND2X1_607 INVX8_10/A OAI21X1_789/Y gnd OAI21X1_790/C vdd NAND2X1
XINVX1_282 NOR2X1_66/A gnd INVX1_282/Y vdd INVX1
XNAND2X1_629 NOR2X1_488/Y OAI22X1_29/Y gnd NOR2X1_489/B vdd NAND2X1
XINVX1_271 BUFX2_21/A gnd INVX1_271/Y vdd INVX1
XNAND2X1_82 XNOR2X1_26/Y XNOR2X1_27/Y gnd NOR2X1_70/A vdd NAND2X1
XNAND2X1_93 MUX2X1_8/S operand_A[25] gnd OAI21X1_44/C vdd NAND2X1
XNAND2X1_60 INVX2_94/A XNOR2X1_46/B gnd NOR2X1_48/A vdd NAND2X1
XNAND2X1_71 XNOR2X1_18/Y XNOR2X1_19/Y gnd OR2X2_3/A vdd NAND2X1
XAOI21X1_231 AOI21X1_231/A OAI21X1_572/Y NOR2X1_326/Y gnd DFFPOSX1_58/D vdd AOI21X1
XAOI21X1_264 INVX1_258/A OAI21X1_600/B OAI21X1_621/B gnd OAI21X1_626/A vdd AOI21X1
XAOI21X1_275 NAND3X1_40/Y AOI21X1_275/B NAND3X1_41/Y gnd AOI21X1_276/B vdd AOI21X1
XAOI21X1_253 INVX4_11/Y OAI21X1_603/Y BUFX4_8/Y gnd OAI22X1_38/A vdd AOI21X1
XAOI21X1_220 INVX1_228/A INVX1_234/Y BUFX4_9/Y gnd OAI22X1_34/A vdd AOI21X1
XAOI21X1_242 BUFX4_167/Y AND2X2_20/Y INVX1_228/Y gnd OAI22X1_18/C vdd AOI21X1
XAOI21X1_286 OAI21X1_653/Y NOR2X1_121/Y OAI21X1_654/Y gnd NAND3X1_54/B vdd AOI21X1
XAOI21X1_297 MUX2X1_5/S operand_A[1] INVX2_58/A gnd AOI21X1_298/B vdd AOI21X1
XOAI21X1_409 INVX2_74/A OAI21X1_409/B OAI21X1_409/C gnd OAI21X1_409/Y vdd OAI21X1
XFILL_21_2 gnd vdd FILL
XFILL_14_1 gnd vdd FILL
XNAND2X1_437 INVX1_157/A INVX1_126/A gnd AND2X2_27/B vdd NAND2X1
XNAND2X1_426 INVX1_190/Y INVX1_191/Y gnd NAND2X1_427/B vdd NAND2X1
XNAND2X1_404 MUX2X1_4/S operand_A[43] gnd OAI21X1_432/C vdd NAND2X1
XNAND2X1_459 NAND2X1_459/A OAI21X1_516/Y gnd NAND2X1_459/Y vdd NAND2X1
XNAND2X1_415 BUFX4_120/Y OAI21X1_441/Y gnd OAI21X1_442/C vdd NAND2X1
XNAND2X1_448 BUFX4_164/Y OAI21X1_234/Y gnd OAI21X1_871/A vdd NAND2X1
XFILL_25_4_1 gnd vdd FILL
XNOR2X1_492 NOR2X1_492/A NOR2X1_492/B gnd NOR2X1_492/Y vdd NOR2X1
XFILL_0_4_1 gnd vdd FILL
XNOR2X1_470 OR2X2_13/B NOR2X1_470/B gnd NOR2X1_470/Y vdd NOR2X1
XNOR2X1_481 XNOR2X1_25/Y INVX1_315/Y gnd OR2X2_46/A vdd NOR2X1
XOAI21X1_943 NOR2X1_3/A NOR2X1_508/Y OAI21X1_943/C gnd OAI21X1_943/Y vdd OAI21X1
XOAI21X1_932 operand_B[26] INVX2_31/Y OAI21X1_932/C gnd XNOR2X1_48/A vdd OAI21X1
XOAI21X1_921 OAI21X1_23/A OR2X2_2/B OAI21X1_22/B gnd INVX1_325/A vdd OAI21X1
XOAI21X1_910 OAI21X1_34/A NAND2X1_59/B BUFX4_141/Y gnd OAI21X1_910/Y vdd OAI21X1
XINVX2_51 operand_B[31] gnd INVX2_51/Y vdd INVX2
XINVX2_40 operand_A[52] gnd INVX2_40/Y vdd INVX2
XINVX2_62 INVX2_62/A gnd INVX2_62/Y vdd INVX2
XINVX2_73 operand_A[43] gnd INVX2_73/Y vdd INVX2
XFILL_7_0_0 gnd vdd FILL
XFILL_8_5_1 gnd vdd FILL
XINVX2_84 INVX2_84/A gnd INVX2_84/Y vdd INVX2
XFILL_16_4_1 gnd vdd FILL
XOAI21X1_25 operand_B[28] INVX4_2/Y NAND2X1_3/A gnd AND2X2_2/A vdd OAI21X1
XOAI21X1_47 INVX2_35/Y MUX2X1_5/S OAI21X1_47/C gnd OAI21X1_47/Y vdd OAI21X1
XOAI21X1_69 BUFX4_68/Y OAI21X1_69/B OAI21X1_69/C gnd OAI21X1_73/A vdd OAI21X1
XOAI21X1_58 MUX2X1_98/S MUX2X1_4/Y OAI21X1_58/C gnd OAI21X1_58/Y vdd OAI21X1
XOAI21X1_14 NOR2X1_24/A OAI21X1_14/B AOI21X1_8/Y gnd AOI21X1_9/C vdd OAI21X1
XOAI21X1_36 INVX2_6/Y BUFX4_46/Y OAI21X1_36/C gnd INVX1_36/A vdd OAI21X1
XOAI21X1_239 INVX4_16/A INVX4_15/A OAI21X1_239/C gnd INVX1_108/A vdd OAI21X1
XOAI21X1_217 INVX2_56/Y MUX2X1_8/S OAI21X1_217/C gnd INVX1_105/A vdd OAI21X1
XOAI21X1_206 INVX8_8/Y NAND3X1_7/Y INVX8_15/Y gnd OAI21X1_222/C vdd OAI21X1
XOAI21X1_228 OAI21X1_228/A BUFX4_22/Y OAI21X1_228/C gnd OR2X2_7/A vdd OAI21X1
XAND2X2_28 AND2X2_28/A AND2X2_28/B gnd AND2X2_28/Y vdd AND2X2
XAND2X2_17 INVX1_163/Y AND2X2_17/B gnd AND2X2_17/Y vdd AND2X2
XAND2X2_39 AND2X2_39/A AND2X2_39/B gnd AND2X2_40/B vdd AND2X2
XNAND2X1_212 BUFX4_36/Y OAI21X1_178/Y gnd OAI21X1_179/C vdd NAND2X1
XNAND2X1_234 BUFX4_18/Y OAI21X1_374/B gnd OAI21X1_201/C vdd NAND2X1
XNAND2X1_223 BUFX4_74/Y OAI21X1_54/B gnd OAI21X1_190/C vdd NAND2X1
XNAND2X1_201 operand_A[9] INVX2_25/Y gnd OAI21X1_639/C vdd NAND2X1
XNAND2X1_267 operand_A[34] operand_B[34] gnd INVX4_17/A vdd NAND2X1
XNAND2X1_289 OAI21X1_283/C AOI22X1_6/D gnd INVX2_62/A vdd NAND2X1
XNAND2X1_256 BUFX4_72/Y INVX1_71/A gnd OAI21X1_227/C vdd NAND2X1
XNAND2X1_278 BUFX4_119/Y INVX1_37/A gnd OAI21X1_254/C vdd NAND2X1
XNAND2X1_245 BUFX4_179/Y OAI21X1_213/Y gnd OAI21X1_221/C vdd NAND2X1
XOAI21X1_784 BUFX4_131/Y INVX1_295/A OAI21X1_784/C gnd MUX2X1_122/A vdd OAI21X1
XOAI21X1_773 INVX1_302/A XNOR2X1_19/Y BUFX4_140/Y gnd OAI21X1_777/B vdd OAI21X1
XOAI21X1_751 OAI21X1_9/Y NAND3X1_4/B BUFX4_105/Y gnd NOR2X1_439/A vdd OAI21X1
XOAI21X1_795 INVX1_305/Y BUFX4_62/Y OAI21X1_795/C gnd OR2X2_42/A vdd OAI21X1
XOAI21X1_740 MUX2X1_102/Y OR2X2_7/B AND2X2_11/B gnd OAI21X1_740/Y vdd OAI21X1
XOAI21X1_762 BUFX4_125/Y OAI21X1_762/B OAI21X1_762/C gnd NOR2X1_471/B vdd OAI21X1
XFILL_31_2_1 gnd vdd FILL
XBUFX4_80 INVX8_4/Y gnd BUFX4_80/Y vdd BUFX4
XBUFX4_91 BUFX4_91/A gnd BUFX4_91/Y vdd BUFX4
XFILL_22_2_1 gnd vdd FILL
XXNOR2X1_1 operand_A[30] operand_B[30] gnd INVX4_1/A vdd XNOR2X1
XFILL_5_3_1 gnd vdd FILL
XINVX1_1 operand_B[28] gnd INVX1_1/Y vdd INVX1
XFILL_13_2_1 gnd vdd FILL
XOAI21X1_592 INVX1_238/Y BUFX4_70/Y OAI21X1_592/C gnd OAI21X1_630/A vdd OAI21X1
XOAI21X1_581 OAI21X1_581/A INVX8_4/A OAI21X1_581/C gnd OAI21X1_581/Y vdd OAI21X1
XOAI21X1_570 OAI22X1_1/B OR2X2_43/A OAI21X1_570/C gnd OAI22X1_34/D vdd OAI21X1
XINVX4_19 INVX4_19/A gnd INVX4_19/Y vdd INVX4
XAND2X2_1 NOR2X1_6/Y AND2X2_1/B gnd AND2X2_1/Y vdd AND2X2
XFILL_2_1 gnd vdd FILL
XAOI21X1_413 BUFX4_141/Y XNOR2X1_49/Y OAI21X1_950/Y gnd AOI21X1_414/B vdd AOI21X1
XAOI21X1_402 NOR2X1_67/B INVX1_325/A BUFX4_29/Y gnd OAI21X1_922/C vdd AOI21X1
XNAND3X1_39 BUFX4_107/Y NAND3X1_39/B NAND3X1_39/C gnd NAND3X1_39/Y vdd NAND3X1
XNAND3X1_28 NAND3X1_28/A NAND3X1_28/B INVX8_13/Y gnd NAND3X1_28/Y vdd NAND3X1
XNAND3X1_17 NAND3X1_17/A NAND3X1_17/B NAND3X1_17/C gnd NOR2X1_186/A vdd NAND3X1
XNOR2X1_17 NOR2X1_19/B INVX2_12/Y gnd NOR2X1_17/Y vdd NOR2X1
XNOR2X1_28 XNOR2X1_6/Y XNOR2X1_7/Y gnd NOR2X1_28/Y vdd NOR2X1
XFILL_27_1_1 gnd vdd FILL
XNOR2X1_39 INVX2_15/Y INVX1_15/Y gnd NOR2X1_39/Y vdd NOR2X1
XFILL_2_1_1 gnd vdd FILL
XFILL_10_0_1 gnd vdd FILL
XMUX2X1_68 operand_A[29] operand_A[28] MUX2X1_9/S gnd MUX2X1_69/A vdd MUX2X1
XMUX2X1_13 operand_A[60] operand_A[59] MUX2X1_3/S gnd MUX2X1_13/Y vdd MUX2X1
XMUX2X1_79 operand_A[24] operand_A[23] MUX2X1_7/S gnd MUX2X1_79/Y vdd MUX2X1
XMUX2X1_24 MUX2X1_24/A MUX2X1_24/B MUX2X1_71/S gnd MUX2X1_24/Y vdd MUX2X1
XFILL_18_1_1 gnd vdd FILL
XMUX2X1_57 MUX2X1_57/A MUX2X1_57/B MUX2X1_57/S gnd MUX2X1_57/Y vdd MUX2X1
XNOR2X1_129 BUFX4_83/Y INVX8_7/Y gnd INVX4_18/A vdd NOR2X1
XMUX2X1_35 MUX2X1_35/A MUX2X1_35/B MUX2X1_2/S gnd MUX2X1_35/Y vdd MUX2X1
XNOR2X1_118 operand_A[11] INVX2_28/Y gnd NOR2X1_118/Y vdd NOR2X1
XNOR2X1_107 XNOR2X1_16/Y XNOR2X1_17/Y gnd NOR2X1_107/Y vdd NOR2X1
XMUX2X1_46 MUX2X1_46/A MUX2X1_46/B MUX2X1_49/S gnd MUX2X1_46/Y vdd MUX2X1
XINVX1_250 INVX1_250/A gnd INVX1_250/Y vdd INVX1
XINVX1_261 INVX1_261/A gnd INVX1_261/Y vdd INVX1
XINVX1_283 INVX1_283/A gnd INVX1_283/Y vdd INVX1
XNAND2X1_50 OAI21X1_33/C NAND2X1_50/B gnd NOR2X1_67/B vdd NAND2X1
XINVX1_294 MUX2X1_78/Y gnd INVX1_294/Y vdd INVX1
XNAND2X1_61 AND2X2_71/B XNOR2X1_13/Y gnd NOR2X1_48/B vdd NAND2X1
XNAND2X1_608 NAND2X1_608/A NOR2X1_451/Y gnd OAI21X1_791/A vdd NAND2X1
XNAND2X1_619 NAND2X1_619/A OAI21X1_830/Y gnd NAND2X1_619/Y vdd NAND2X1
XINVX1_272 BUFX2_20/A gnd INVX1_272/Y vdd INVX1
XNAND2X1_83 XNOR2X1_47/B XNOR2X1_29/Y gnd NOR2X1_70/B vdd NAND2X1
XNAND2X1_94 BUFX4_69/Y INVX1_95/A gnd OAI21X1_45/C vdd NAND2X1
XNAND2X1_72 XNOR2X1_20/Y XNOR2X1_21/Y gnd OR2X2_3/B vdd NAND2X1
XAOI21X1_210 OR2X2_33/B OAI21X1_552/B BUFX4_32/Y gnd OAI21X1_552/C vdd AOI21X1
XAOI21X1_287 NOR2X1_417/Y INVX2_86/Y NOR2X1_416/Y gnd OAI21X1_658/C vdd AOI21X1
XAOI21X1_276 NAND3X1_39/Y AOI21X1_276/B NOR2X1_375/Y gnd DFFPOSX1_64/D vdd AOI21X1
XAOI21X1_265 OAI21X1_597/C OAI21X1_599/Y INVX1_258/Y gnd OAI21X1_621/A vdd AOI21X1
XAOI21X1_232 NOR2X1_321/A INVX2_82/A NOR2X1_320/B gnd INVX1_246/A vdd AOI21X1
XAOI21X1_254 BUFX4_167/Y MUX2X1_61/Y INVX8_7/Y gnd AOI21X1_255/B vdd AOI21X1
XAOI21X1_221 INVX8_10/A INVX1_234/A OAI22X1_34/A gnd NAND2X1_494/A vdd AOI21X1
XAOI21X1_243 AOI21X1_243/A NAND2X1_508/Y OAI22X1_18/Y gnd OAI21X1_595/A vdd AOI21X1
XAOI21X1_298 BUFX4_66/Y AOI21X1_298/B OAI21X1_692/Y gnd OAI21X1_693/B vdd AOI21X1
XNAND2X1_427 INVX1_194/A NAND2X1_427/B gnd INVX4_22/A vdd NAND2X1
XNAND2X1_405 BUFX4_73/Y OAI21X1_457/B gnd OAI21X1_433/C vdd NAND2X1
XNAND2X1_416 BUFX4_19/Y INVX1_181/Y gnd OAI21X1_443/C vdd NAND2X1
XNAND2X1_449 AND2X2_26/B INVX1_204/A gnd INVX1_207/A vdd NAND2X1
XNAND2X1_438 operand_A[47] INVX1_191/Y gnd OAI21X1_668/C vdd NAND2X1
XOAI21X1_900 AND2X2_73/A INVX2_94/Y BUFX4_108/Y gnd NOR2X1_496/A vdd OAI21X1
XNOR2X1_493 BUFX4_10/Y NOR2X1_493/B gnd OAI22X1_31/C vdd NOR2X1
XNOR2X1_460 NOR2X1_460/A NOR2X1_460/B gnd NOR2X1_460/Y vdd NOR2X1
XNOR2X1_471 OR2X2_39/B NOR2X1_471/B gnd NOR2X1_471/Y vdd NOR2X1
XNOR2X1_482 BUFX4_31/Y OR2X2_46/A gnd NOR2X1_482/Y vdd NOR2X1
XOAI21X1_944 operand_B[28] INVX4_2/Y OAI21X1_944/C gnd XNOR2X1_49/A vdd OAI21X1
XOAI21X1_922 NOR2X1_67/B INVX1_325/A OAI21X1_922/C gnd AOI22X1_56/D vdd OAI21X1
XOAI21X1_911 INVX1_234/Y BUFX4_171/Y BUFX4_114/Y gnd OAI22X1_34/B vdd OAI21X1
XOAI21X1_933 OAI22X1_18/B INVX2_49/Y NOR2X1_22/A gnd OAI22X1_37/B vdd OAI21X1
XINVX2_63 INVX2_63/A gnd INVX2_63/Y vdd INVX2
XINVX2_52 operand_A[49] gnd INVX2_52/Y vdd INVX2
XINVX2_41 operand_A[50] gnd INVX2_41/Y vdd INVX2
XINVX2_85 operand_A[59] gnd INVX2_85/Y vdd INVX2
XINVX2_74 INVX2_74/A gnd OR2X2_21/B vdd INVX2
XINVX2_30 operand_A[27] gnd INVX2_30/Y vdd INVX2
XFILL_7_0_1 gnd vdd FILL
XOAI21X1_48 INVX1_41/Y BUFX4_69/Y OAI21X1_48/C gnd OAI21X1_48/Y vdd OAI21X1
XOAI21X1_15 INVX2_19/Y INVX2_18/Y NAND3X1_1/A gnd NOR2X1_29/B vdd OAI21X1
XOAI21X1_59 INVX1_45/Y MUX2X1_51/S OAI21X1_59/C gnd INVX1_46/A vdd OAI21X1
XOAI21X1_37 INVX4_5/Y BUFX4_48/Y OAI21X1_37/C gnd INVX1_91/A vdd OAI21X1
XOAI21X1_26 NOR2X1_66/A INVX1_316/A OAI21X1_26/C gnd OAI21X1_26/Y vdd OAI21X1
XAND2X2_29 AND2X2_29/A AND2X2_29/B gnd AND2X2_30/B vdd AND2X2
XOAI21X1_218 INVX1_105/Y MUX2X1_23/S OAI21X1_218/C gnd INVX1_106/A vdd OAI21X1
XOAI21X1_229 BUFX4_192/Y OAI21X1_229/B OAI21X1_229/C gnd OAI21X1_231/B vdd OAI21X1
XAND2X2_18 AND2X2_18/A NOR2X1_80/A gnd AND2X2_18/Y vdd AND2X2
XOAI21X1_207 XOR2X1_3/A INVX1_68/A OAI21X1_207/C gnd MUX2X1_35/A vdd OAI21X1
XNAND2X1_268 AOI22X1_4/C INVX4_16/Y gnd OAI21X1_240/B vdd NAND2X1
XNAND2X1_213 BUFX4_71/Y OAI21X1_76/B gnd OAI21X1_180/C vdd NAND2X1
XNAND2X1_202 operand_A[8] INVX1_20/Y gnd OAI21X1_806/C vdd NAND2X1
XNAND2X1_224 BUFX4_74/Y OAI21X1_57/Y gnd OAI21X1_191/C vdd NAND2X1
XNAND2X1_246 BUFX4_191/Y OAI21X1_99/Y gnd OAI21X1_214/C vdd NAND2X1
XNAND2X1_235 BUFX4_162/Y NOR2X1_128/Y gnd INVX1_100/A vdd NAND2X1
XNAND2X1_257 BUFX4_22/Y MUX2X1_27/Y gnd OAI21X1_228/C vdd NAND2X1
XNAND2X1_279 BUFX4_17/Y INVX1_112/Y gnd OAI21X1_255/C vdd NAND2X1
XNOR2X1_290 operand_A[54] operand_B[54] gnd OAI22X1_13/D vdd NOR2X1
XOAI21X1_741 NOR2X1_19/B INVX2_12/Y OAI21X1_741/C gnd OAI21X1_742/B vdd OAI21X1
XOAI21X1_730 NOR2X1_428/A NOR2X1_15/Y XOR2X1_7/Y gnd OAI21X1_741/C vdd OAI21X1
XOAI21X1_752 XNOR2X1_21/Y OAI21X1_28/Y OAI21X1_752/C gnd OAI21X1_752/Y vdd OAI21X1
XOAI21X1_774 operand_A[6] operand_B[6] BUFX4_2/Y gnd OAI21X1_775/C vdd OAI21X1
XOAI21X1_763 INVX1_299/Y BUFX4_24/Y OAI21X1_763/C gnd NOR2X1_442/B vdd OAI21X1
XOAI21X1_796 BUFX4_41/Y OAI21X1_796/B OAI21X1_796/C gnd OAI21X1_796/Y vdd OAI21X1
XOAI21X1_785 MUX2X1_57/S MUX2X1_115/Y NOR2X1_450/Y gnd OAI21X1_789/C vdd OAI21X1
XBUFX4_70 INVX8_1/Y gnd BUFX4_70/Y vdd BUFX4
XBUFX4_81 INVX8_4/Y gnd BUFX4_81/Y vdd BUFX4
XBUFX4_92 INVX8_11/Y gnd BUFX4_92/Y vdd BUFX4
XOR2X2_40 OR2X2_40/A OR2X2_40/B gnd OR2X2_40/Y vdd OR2X2
XXNOR2X1_2 operand_B[29] operand_A[29] gnd NOR2X1_3/A vdd XNOR2X1
XOAI21X1_582 INVX1_232/A INVX1_239/Y INVX1_246/A gnd OAI21X1_583/B vdd OAI21X1
XINVX1_2 INVX1_2/A gnd INVX1_2/Y vdd INVX1
XOAI21X1_571 operand_A[56] operand_B[56] BUFX4_4/Y gnd AND2X2_37/B vdd OAI21X1
XOAI21X1_593 INVX1_227/Y MUX2X1_62/S OAI21X1_593/C gnd MUX2X1_58/A vdd OAI21X1
XOAI21X1_560 OAI21X1_560/A MUX2X1_34/S BUFX4_79/Y gnd NOR2X1_301/B vdd OAI21X1
XFILL_32_5_0 gnd vdd FILL
XFILL_23_5_0 gnd vdd FILL
XFILL_14_5_0 gnd vdd FILL
XAND2X2_2 AND2X2_2/A AND2X2_2/B gnd AND2X2_2/Y vdd AND2X2
XOAI21X1_390 INVX1_167/Y BUFX4_22/Y OAI21X1_390/C gnd AND2X2_18/A vdd OAI21X1
XAOI21X1_414 OAI21X1_943/Y AOI21X1_414/B NOR2X1_511/Y gnd DFFPOSX1_30/D vdd AOI21X1
XAOI21X1_403 XNOR2X1_27/Y OAI21X1_924/A OAI21X1_924/Y gnd NOR2X1_501/A vdd AOI21X1
XNAND3X1_29 OR2X2_28/Y NAND3X1_29/B NAND3X1_29/C gnd NAND3X1_29/Y vdd NAND3X1
XNAND3X1_18 NAND3X1_18/A NAND3X1_18/B NOR2X1_199/Y gnd NAND3X1_18/Y vdd NAND3X1
XNOR2X1_18 NOR2X1_83/A INVX2_12/Y gnd OAI21X1_8/A vdd NOR2X1
XNOR2X1_29 NOR2X1_29/A NOR2X1_29/B gnd NOR2X1_29/Y vdd NOR2X1
XNOR2X1_119 AND2X2_6/Y INVX4_1/Y gnd NOR2X1_119/Y vdd NOR2X1
XMUX2X1_14 operand_A[56] operand_A[55] MUX2X1_8/S gnd MUX2X1_14/Y vdd MUX2X1
XMUX2X1_69 MUX2X1_69/A MUX2X1_7/Y BUFX4_72/Y gnd MUX2X1_71/B vdd MUX2X1
XMUX2X1_36 MUX2X1_36/A MUX2X1_36/B BUFX4_16/Y gnd MUX2X1_36/Y vdd MUX2X1
XMUX2X1_47 MUX2X1_61/A MUX2X1_47/B BUFX4_18/Y gnd MUX2X1_47/Y vdd MUX2X1
XMUX2X1_58 MUX2X1_58/A MUX2X1_58/B BUFX4_18/Y gnd MUX2X1_58/Y vdd MUX2X1
XNOR2X1_108 XNOR2X1_18/Y XNOR2X1_19/Y gnd NAND3X1_4/C vdd NOR2X1
XMUX2X1_25 MUX2X1_42/B MUX2X1_25/B MUX2X1_25/S gnd MUX2X1_25/Y vdd MUX2X1
XINVX1_273 BUFX2_19/A gnd INVX1_273/Y vdd INVX1
XINVX1_240 INVX1_240/A gnd INVX1_240/Y vdd INVX1
XINVX1_251 INVX1_251/A gnd INVX1_251/Y vdd INVX1
XINVX1_284 MUX2X1_73/Y gnd INVX1_284/Y vdd INVX1
XINVX1_262 BUFX2_14/A gnd INVX1_262/Y vdd INVX1
XINVX1_295 INVX1_295/A gnd INVX1_295/Y vdd INVX1
XNAND2X1_609 INVX8_5/A MUX2X1_126/B gnd NAND2X1_609/Y vdd NAND2X1
XNAND2X1_84 NOR2X1_3/A NOR2X1_3/B gnd INVX1_34/A vdd NAND2X1
XNAND2X1_51 NOR2X1_67/A NOR2X1_67/B gnd OR2X2_2/A vdd NAND2X1
XNAND2X1_95 MUX2X1_4/S operand_A[27] gnd OAI21X1_46/C vdd NAND2X1
XNAND2X1_40 XNOR2X1_41/B NAND2X1_40/B gnd NOR2X1_29/A vdd NAND2X1
XNAND2X1_73 BUFX4_113/Y INVX2_14/Y gnd NAND2X1_73/Y vdd NAND2X1
XNAND2X1_62 XNOR2X1_14/Y XNOR2X1_15/Y gnd NOR2X1_66/A vdd NAND2X1
XAOI21X1_200 INVX1_224/A OAI21X1_544/B BUFX4_32/Y gnd OAI21X1_544/C vdd AOI21X1
XAOI21X1_211 OR2X2_33/B OR2X2_33/A BUFX4_93/Y gnd AOI21X1_214/A vdd AOI21X1
XAOI21X1_233 INVX2_84/A OAI21X1_583/B BUFX4_30/Y gnd OAI21X1_583/C vdd AOI21X1
XAOI21X1_288 NOR2X1_310/Y OAI21X1_661/Y OAI21X1_660/Y gnd OAI21X1_662/C vdd AOI21X1
XAOI21X1_266 INVX2_89/Y OAI21X1_610/Y INVX1_260/A gnd OAI21X1_627/A vdd AOI21X1
XFILL_20_3_0 gnd vdd FILL
XAOI21X1_222 BUFX4_80/Y NAND2X1_494/Y NAND3X1_34/Y gnd AND2X2_38/B vdd AOI21X1
XAOI21X1_244 BUFX4_113/Y OAI22X1_37/D OR2X2_35/Y gnd OAI21X1_595/C vdd AOI21X1
XAOI21X1_255 NAND2X1_513/Y AOI21X1_255/B OAI22X1_38/A gnd OAI21X1_607/A vdd AOI21X1
XAOI21X1_277 OAI21X1_8/B XNOR2X1_17/Y INVX1_280/Y gnd OAI21X1_643/C vdd AOI21X1
XAOI21X1_299 INVX2_10/Y BUFX4_150/Y OAI21X1_697/Y gnd AND2X2_51/A vdd AOI21X1
XFILL_28_4_0 gnd vdd FILL
XFILL_3_4_0 gnd vdd FILL
XFILL_11_3_0 gnd vdd FILL
XFILL_19_4_0 gnd vdd FILL
XNAND2X1_439 BUFX4_73/Y OAI21X1_504/B gnd OAI21X1_480/C vdd NAND2X1
XNAND2X1_406 INVX8_3/A OAI21X1_372/Y gnd OAI21X1_434/C vdd NAND2X1
XNAND2X1_417 NAND2X1_417/A NAND2X1_417/B gnd NAND3X1_24/C vdd NAND2X1
XNAND2X1_428 BUFX4_164/Y OAI21X1_123/A gnd INVX1_193/A vdd NAND2X1
XOAI21X1_901 OAI21X1_901/A NOR2X1_48/B OAI21X1_27/B gnd OAI21X1_902/B vdd OAI21X1
XOAI21X1_934 operand_B[27] operand_A[27] BUFX4_6/Y gnd OAI21X1_935/C vdd OAI21X1
XOAI21X1_923 OAI21X1_34/A NOR2X1_70/B INVX1_32/A gnd OAI21X1_924/A vdd OAI21X1
XOAI21X1_912 BUFX4_158/Y NOR2X1_42/Y OAI22X1_3/C gnd OAI21X1_913/C vdd OAI21X1
XNOR2X1_494 INVX8_7/Y OR2X2_32/A gnd OAI22X1_31/A vdd NOR2X1
XNOR2X1_472 XNOR2X1_23/Y NOR2X1_472/B gnd INVX1_313/A vdd NOR2X1
XNOR2X1_461 MUX2X1_64/S NOR2X1_461/B gnd NOR2X1_462/A vdd NOR2X1
XNOR2X1_483 NOR2X1_483/A NOR2X1_483/B gnd AND2X2_67/B vdd NOR2X1
XNOR2X1_450 BUFX4_111/Y NOR2X1_450/B gnd NOR2X1_450/Y vdd NOR2X1
XOAI21X1_945 BUFX4_163/Y OAI21X1_945/B OAI21X1_945/C gnd AOI22X1_58/C vdd OAI21X1
XINVX2_86 OR2X2_34/B gnd INVX2_86/Y vdd INVX2
XINVX2_64 INVX2_64/A gnd INVX2_64/Y vdd INVX2
XINVX2_42 operand_A[48] gnd INVX2_42/Y vdd INVX2
XINVX2_53 operand_A[53] gnd INVX2_53/Y vdd INVX2
XINVX2_75 INVX2_75/A gnd INVX2_75/Y vdd INVX2
XINVX2_31 operand_A[26] gnd INVX2_31/Y vdd INVX2
XINVX2_20 operand_A[13] gnd INVX2_20/Y vdd INVX2
XOAI21X1_16 NOR2X1_30/Y NOR2X1_31/Y XOR2X1_6/Y gnd OAI21X1_17/A vdd OAI21X1
XOAI21X1_27 NOR2X1_48/A OAI21X1_27/B OAI21X1_27/C gnd INVX1_28/A vdd OAI21X1
XOAI21X1_38 INVX1_36/Y BUFX4_67/Y OAI21X1_38/C gnd INVX1_37/A vdd OAI21X1
XOAI21X1_49 INVX1_40/Y BUFX4_119/Y OAI21X1_49/C gnd INVX1_42/A vdd OAI21X1
XOAI21X1_219 INVX1_63/Y XOR2X1_3/A OAI21X1_219/C gnd OAI21X1_219/Y vdd OAI21X1
XOAI21X1_208 INVX1_102/Y BUFX4_76/Y OAI21X1_208/C gnd INVX1_136/A vdd OAI21X1
XAND2X2_19 AND2X2_19/A INVX8_11/A gnd AND2X2_19/Y vdd AND2X2
XNAND2X1_236 operand_A[33] operand_B[33] gnd OAI21X1_239/C vdd NAND2X1
XNAND2X1_214 BUFX4_72/Y OAI21X1_77/Y gnd OAI21X1_181/C vdd NAND2X1
XNAND2X1_258 BUFX4_191/Y MUX2X1_14/Y gnd OAI21X1_229/C vdd NAND2X1
XNAND2X1_269 MUX2X1_30/S INVX1_50/Y gnd OAI21X1_245/C vdd NAND2X1
XNAND2X1_225 MUX2X1_2/S OAI21X1_290/B gnd OAI21X1_192/C vdd NAND2X1
XNAND2X1_203 operand_A[10] INVX2_23/Y gnd OAI21X1_162/B vdd NAND2X1
XNAND2X1_247 MUX2X1_97/S OAI21X1_96/Y gnd OAI21X1_215/C vdd NAND2X1
XFILL_25_2_0 gnd vdd FILL
XFILL_0_2_0 gnd vdd FILL
XNOR2X1_280 BUFX4_32/Y NOR2X1_286/B gnd NOR2X1_280/Y vdd NOR2X1
XNOR2X1_291 OAI22X1_13/D AND2X2_33/Y gnd INVX1_224/A vdd NOR2X1
XOAI21X1_720 MUX2X1_76/A BUFX4_66/Y NOR2X1_19/B gnd OAI21X1_721/B vdd OAI21X1
XOAI21X1_731 XOR2X1_7/A operand_A[2] BUFX4_2/Y gnd NAND3X1_57/B vdd OAI21X1
XOAI21X1_742 XOR2X1_4/Y OAI21X1_742/B OAI21X1_742/C gnd NAND3X1_59/A vdd OAI21X1
XOAI21X1_775 BUFX4_154/Y XNOR2X1_19/Y OAI21X1_775/C gnd OR2X2_41/A vdd OAI21X1
XOAI21X1_753 BUFX4_183/Y operand_A[4] BUFX4_2/Y gnd OAI21X1_754/C vdd OAI21X1
XOAI21X1_764 INVX1_300/Y AND2X2_56/Y BUFX4_90/Y gnd NAND3X1_62/A vdd OAI21X1
XOAI21X1_786 OR2X2_15/A BUFX4_77/Y OAI21X1_789/C gnd OAI21X1_786/Y vdd OAI21X1
XFILL_8_3_0 gnd vdd FILL
XOAI21X1_797 NOR2X1_452/Y OAI21X1_800/B BUFX4_89/Y gnd OAI21X1_797/Y vdd OAI21X1
XFILL_16_2_0 gnd vdd FILL
XBUFX4_93 INVX8_11/Y gnd BUFX4_93/Y vdd BUFX4
XBUFX4_71 INVX8_1/Y gnd BUFX4_71/Y vdd BUFX4
XBUFX4_60 BUFX4_60/A gnd BUFX4_60/Y vdd BUFX4
XBUFX4_82 INVX8_4/Y gnd BUFX4_82/Y vdd BUFX4
XXNOR2X1_3 operand_B[28] operand_A[28] gnd NOR2X1_3/B vdd XNOR2X1
XOR2X2_30 OR2X2_30/A OR2X2_30/B gnd OR2X2_30/Y vdd OR2X2
XOR2X2_41 OR2X2_41/A OR2X2_41/B gnd OR2X2_41/Y vdd OR2X2
XOR2X2_1 OR2X2_1/A OR2X2_1/B gnd OR2X2_1/Y vdd OR2X2
XOAI21X1_583 INVX2_84/A OAI21X1_583/B OAI21X1_583/C gnd OAI21X1_583/Y vdd OAI21X1
XOAI21X1_572 INVX2_82/Y NOR2X1_321/Y OAI21X1_572/C gnd OAI21X1_572/Y vdd OAI21X1
XOAI21X1_594 BUFX4_64/Y INVX1_243/Y AOI22X1_27/Y gnd OR2X2_35/A vdd OAI21X1
XOAI21X1_550 OAI21X1_903/A BUFX4_174/Y AND2X2_34/Y gnd OAI21X1_550/Y vdd OAI21X1
XINVX1_3 INVX1_3/A gnd INVX1_3/Y vdd INVX1
XOAI21X1_561 NOR2X1_301/Y NOR2X1_299/Y INVX8_7/A gnd OAI21X1_561/Y vdd OAI21X1
XFILL_32_5_1 gnd vdd FILL
XFILL_31_0_0 gnd vdd FILL
XFILL_23_5_1 gnd vdd FILL
XFILL_22_0_0 gnd vdd FILL
XFILL_5_1_0 gnd vdd FILL
XFILL_14_5_1 gnd vdd FILL
XFILL_13_0_0 gnd vdd FILL
XOAI21X1_380 INVX1_163/A INVX1_154/A AND2X2_16/Y gnd OAI21X1_380/Y vdd OAI21X1
XAND2X2_3 AND2X2_3/A INVX8_12/A gnd AND2X2_3/Y vdd AND2X2
XOAI21X1_391 INVX1_168/Y OR2X2_13/B INVX2_48/Y gnd OAI21X1_391/Y vdd OAI21X1
XAOI21X1_404 BUFX4_81/Y OAI21X1_925/Y INVX8_9/Y gnd OAI22X1_36/C vdd AOI21X1
XNAND3X1_19 NAND3X1_19/A OR2X2_19/Y NAND3X1_19/C gnd NAND3X1_19/Y vdd NAND3X1
XNOR2X1_19 operand_A[2] NOR2X1_19/B gnd OAI21X1_8/B vdd NOR2X1
XMUX2X1_15 operand_A[48] operand_A[47] MUX2X1_9/S gnd MUX2X1_15/Y vdd MUX2X1
XMUX2X1_59 MUX2X1_65/B MUX2X1_59/B BUFX4_75/Y gnd MUX2X1_60/A vdd MUX2X1
XMUX2X1_48 MUX2X1_48/A MUX2X1_48/B BUFX4_81/Y gnd MUX2X1_48/Y vdd MUX2X1
XMUX2X1_37 MUX2X1_43/B MUX2X1_37/B BUFX4_25/Y gnd MUX2X1_37/Y vdd MUX2X1
XNOR2X1_109 OR2X2_1/A OR2X2_1/B gnd NOR2X1_109/Y vdd NOR2X1
XMUX2X1_26 MUX2X1_37/B MUX2X1_26/B BUFX4_23/Y gnd MUX2X1_44/B vdd MUX2X1
XINVX1_241 INVX1_241/A gnd INVX1_241/Y vdd INVX1
XINVX1_230 operand_B[56] gnd INVX1_230/Y vdd INVX1
XINVX1_252 operand_B[61] gnd INVX1_252/Y vdd INVX1
XINVX1_274 BUFX2_30/A gnd INVX1_274/Y vdd INVX1
XINVX1_296 INVX1_296/A gnd INVX1_296/Y vdd INVX1
XINVX1_285 INVX1_285/A gnd INVX1_285/Y vdd INVX1
XINVX1_263 BUFX2_13/A gnd INVX1_263/Y vdd INVX1
XNAND2X1_96 BUFX4_46/Y operand_A[29] gnd OAI21X1_47/C vdd NAND2X1
XNAND2X1_52 INVX4_8/Y INVX1_23/Y gnd NAND2X1_52/Y vdd NAND2X1
XNAND2X1_30 INVX1_30/A INVX1_85/A gnd NAND3X1_1/A vdd NAND2X1
XNAND2X1_85 MUX2X1_9/S operand_A[15] gnd OAI21X1_36/C vdd NAND2X1
XNAND2X1_74 XNOR2X1_22/Y XNOR2X1_23/Y gnd NOR2X1_59/A vdd NAND2X1
XNAND2X1_41 INVX2_24/Y INVX2_25/Y gnd NAND2X1_41/Y vdd NAND2X1
XNAND2X1_63 operand_B[19] INVX2_7/Y gnd NAND2X1_63/Y vdd NAND2X1
XAOI21X1_223 OAI21X1_564/Y AND2X2_38/Y NOR2X1_303/Y gnd DFFPOSX1_57/D vdd AOI21X1
XAOI21X1_201 NOR2X1_292/Y OAI21X1_532/C OAI21X1_546/Y gnd INVX1_225/A vdd AOI21X1
XFILL_20_3_1 gnd vdd FILL
XAOI21X1_234 INVX4_11/Y NAND2X1_503/Y BUFX4_8/Y gnd OAI22X1_36/A vdd AOI21X1
XAOI21X1_212 BUFX4_163/Y NOR2X1_177/Y INVX1_228/Y gnd OAI22X1_14/C vdd AOI21X1
XAOI21X1_245 AOI21X1_245/A OR2X2_34/Y OAI21X1_595/Y gnd AOI21X1_246/B vdd AOI21X1
XAOI21X1_267 INVX1_259/A OAI21X1_627/A BUFX4_94/Y gnd AOI21X1_271/A vdd AOI21X1
XAOI21X1_289 OAI21X1_656/Y OAI21X1_663/Y OR2X2_38/B gnd NOR2X1_424/A vdd AOI21X1
XAOI21X1_256 INVX4_18/A AND2X2_75/A OAI21X1_606/Y gnd OAI21X1_607/C vdd AOI21X1
XAOI22X1_50 INVX8_7/A MUX2X1_48/B AOI22X1_50/C INVX8_9/A gnd AOI22X1_50/Y vdd AOI22X1
XAOI21X1_278 OAI21X1_158/C INVX2_92/Y NOR2X1_23/Y gnd OAI21X1_644/A vdd AOI21X1
XFILL_28_4_1 gnd vdd FILL
XFILL_3_4_1 gnd vdd FILL
XFILL_11_3_1 gnd vdd FILL
XOAI22X1_1 OAI22X1_1/A OAI22X1_1/B OAI22X1_1/C INVX8_8/Y gnd OAI22X1_2/D vdd OAI22X1
XFILL_19_4_1 gnd vdd FILL
XNAND2X1_407 operand_A[45] operand_B[45] gnd INVX1_182/A vdd NAND2X1
XNAND2X1_429 BUFX4_73/Y OAI21X1_467/Y gnd OAI21X1_468/C vdd NAND2X1
XNAND2X1_418 BUFX4_36/Y NOR2X1_166/B gnd OAI21X1_444/C vdd NAND2X1
XNOR2X1_440 NOR2X1_440/A NOR2X1_440/B gnd NOR2X1_440/Y vdd NOR2X1
XNOR2X1_451 NOR2X1_451/A NOR2X1_451/B gnd NOR2X1_451/Y vdd NOR2X1
XOAI21X1_924 OAI21X1_924/A XNOR2X1_27/Y BUFX4_141/Y gnd OAI21X1_924/Y vdd OAI21X1
XOAI21X1_935 BUFX4_63/Y OAI21X1_935/B OAI21X1_935/C gnd NOR2X1_503/B vdd OAI21X1
XOAI21X1_913 operand_A[24] operand_B[24] OAI21X1_913/C gnd NAND3X1_72/A vdd OAI21X1
XOAI21X1_946 OAI21X1_946/A BUFX4_169/Y BUFX4_112/Y gnd NOR2X1_509/B vdd OAI21X1
XNOR2X1_473 BUFX4_83/Y OR2X2_25/A gnd NOR2X1_473/Y vdd NOR2X1
XNOR2X1_495 NOR2X1_495/A NOR2X1_495/B gnd NOR2X1_495/Y vdd NOR2X1
XOAI21X1_902 INVX2_94/A OAI21X1_902/B OAI21X1_902/C gnd OAI21X1_902/Y vdd OAI21X1
XNOR2X1_462 NOR2X1_462/A NOR2X1_462/B gnd NOR2X1_462/Y vdd NOR2X1
XNOR2X1_484 INVX8_7/Y NOR2X1_484/B gnd OAI22X1_28/D vdd NOR2X1
XINVX2_21 operand_A[12] gnd INVX2_21/Y vdd INVX2
XINVX2_10 INVX2_10/A gnd INVX2_10/Y vdd INVX2
XINVX2_76 operand_B[50] gnd INVX2_76/Y vdd INVX2
XINVX2_65 INVX2_65/A gnd INVX2_65/Y vdd INVX2
XINVX2_54 operand_A[41] gnd INVX2_54/Y vdd INVX2
XINVX2_87 operand_A[60] gnd INVX2_87/Y vdd INVX2
XINVX2_43 operand_A[46] gnd INVX2_43/Y vdd INVX2
XINVX2_32 operand_A[24] gnd INVX2_32/Y vdd INVX2
XOAI21X1_28 OAI21X1_28/A OAI21X1_28/B OAI21X1_28/C gnd OAI21X1_28/Y vdd OAI21X1
XOAI21X1_17 OAI21X1_17/A OAI21X1_17/B OAI21X1_17/C gnd OAI21X1_17/Y vdd OAI21X1
XOAI21X1_39 INVX2_4/Y BUFX4_50/Y OAI21X1_39/C gnd INVX1_38/A vdd OAI21X1
XOAI21X1_209 BUFX4_134/Y INVX1_136/A OAI21X1_209/C gnd OAI21X1_213/B vdd OAI21X1
XFILL_12_1 gnd vdd FILL
XNAND2X1_204 INVX1_34/Y NOR2X1_119/Y gnd NOR2X1_120/A vdd NAND2X1
XNAND2X1_237 OAI21X1_239/C OR2X2_6/Y gnd INVX4_16/A vdd NAND2X1
XNAND2X1_259 BUFX4_71/Y OAI21X1_129/Y gnd OAI21X1_230/C vdd NAND2X1
XNAND2X1_215 BUFX4_71/Y OAI21X1_80/Y gnd OAI21X1_182/C vdd NAND2X1
XNAND2X1_248 MUX2X1_87/S OAI21X1_215/Y gnd OAI21X1_216/C vdd NAND2X1
XNAND2X1_226 OR2X2_13/B OAI21X1_369/A gnd OAI21X1_193/C vdd NAND2X1
XNOR2X1_292 INVX2_78/A INVX1_219/A gnd NOR2X1_292/Y vdd NOR2X1
XNOR2X1_281 INVX4_23/A INVX1_212/A gnd NOR2X1_281/Y vdd NOR2X1
XNOR2X1_270 INVX1_211/Y INVX2_77/Y gnd NOR2X1_271/B vdd NOR2X1
XFILL_25_2_1 gnd vdd FILL
XFILL_0_2_1 gnd vdd FILL
XOAI21X1_798 operand_A[8] operand_B[8] BUFX4_2/Y gnd OAI21X1_799/C vdd OAI21X1
XOAI21X1_787 operand_B[7] operand_A[7] BUFX4_2/Y gnd OAI21X1_788/C vdd OAI21X1
XOAI21X1_743 OAI21X1_28/B OAI21X1_8/B OAI21X1_743/C gnd OAI21X1_744/B vdd OAI21X1
XOAI21X1_721 NOR2X1_432/Y OAI21X1_721/B OAI21X1_721/C gnd MUX2X1_96/B vdd OAI21X1
XOAI21X1_776 BUFX4_62/Y INVX1_303/Y BUFX4_97/Y gnd OR2X2_41/B vdd OAI21X1
XOAI21X1_754 BUFX4_154/Y XNOR2X1_21/Y OAI21X1_754/C gnd NOR2X1_440/B vdd OAI21X1
XOAI21X1_710 MUX2X1_98/S OAI21X1_710/B OAI21X1_710/C gnd INVX1_290/A vdd OAI21X1
XOAI21X1_765 MUX2X1_34/Y BUFX4_82/Y OR2X2_40/Y gnd OAI21X1_765/Y vdd OAI21X1
XOAI21X1_732 NOR2X1_435/Y AND2X2_54/Y BUFX4_112/Y gnd OAI21X1_732/Y vdd OAI21X1
XFILL_8_3_1 gnd vdd FILL
XFILL_16_2_1 gnd vdd FILL
XBUFX4_61 INVX8_17/Y gnd BUFX4_61/Y vdd BUFX4
XBUFX4_50 operand_B[0] gnd BUFX4_50/Y vdd BUFX4
XBUFX4_94 INVX8_11/Y gnd BUFX4_94/Y vdd BUFX4
XBUFX4_72 INVX8_1/Y gnd BUFX4_72/Y vdd BUFX4
XBUFX4_83 INVX8_4/Y gnd BUFX4_83/Y vdd BUFX4
XOR2X2_2 OR2X2_2/A OR2X2_2/B gnd OR2X2_2/Y vdd OR2X2
XOR2X2_20 OR2X2_20/A OR2X2_8/B gnd OR2X2_20/Y vdd OR2X2
XOR2X2_31 OR2X2_31/A OR2X2_31/B gnd OR2X2_31/Y vdd OR2X2
XXNOR2X1_4 operand_A[13] operand_B[13] gnd XNOR2X1_4/Y vdd XNOR2X1
XOR2X2_42 OR2X2_42/A OR2X2_42/B gnd OR2X2_42/Y vdd OR2X2
XINVX1_4 INVX1_4/A gnd INVX1_4/Y vdd INVX1
XOAI21X1_573 OAI21X1_610/A INVX2_81/A NOR2X1_323/Y gnd OAI21X1_573/Y vdd OAI21X1
XOAI21X1_584 INVX4_13/Y operand_B[57] OAI21X1_584/C gnd INVX1_240/A vdd OAI21X1
XOAI21X1_595 OAI21X1_595/A BUFX4_114/Y OAI21X1_595/C gnd OAI21X1_595/Y vdd OAI21X1
XOAI21X1_551 OAI21X1_551/A OR2X2_40/B OAI21X1_551/C gnd OAI21X1_551/Y vdd OAI21X1
XOAI21X1_562 OR2X2_7/B BUFX4_38/Y operand_A[63] gnd INVX1_228/A vdd OAI21X1
XOAI21X1_540 NOR2X1_166/B INVX8_2/A NOR2X1_75/A gnd OAI21X1_541/C vdd OAI21X1
XNAND2X1_590 NOR2X1_54/A OAI21X1_704/Y gnd OAI21X1_735/C vdd NAND2X1
XFILL_31_0_1 gnd vdd FILL
XFILL_22_0_1 gnd vdd FILL
XFILL_5_1_1 gnd vdd FILL
XFILL_13_0_1 gnd vdd FILL
XOAI21X1_381 INVX1_162/A AND2X2_16/B INVX8_11/A gnd NOR2X1_192/A vdd OAI21X1
XAND2X2_4 AND2X2_4/A BUFX4_99/Y gnd AND2X2_4/Y vdd AND2X2
XOAI21X1_392 INVX1_155/Y NOR2X1_219/A OAI21X1_424/A gnd OAI21X1_393/B vdd OAI21X1
XOAI21X1_370 OR2X2_43/A INVX8_8/Y INVX8_15/Y gnd OAI21X1_377/C vdd OAI21X1
XAOI21X1_405 NOR2X1_67/A OAI21X1_931/B BUFX4_29/Y gnd OAI21X1_931/C vdd AOI21X1
XMUX2X1_16 operand_A[52] operand_A[51] BUFX4_48/Y gnd MUX2X1_16/Y vdd MUX2X1
XMUX2X1_27 MUX2X1_27/A MUX2X1_27/B MUX2X1_27/S gnd MUX2X1_27/Y vdd MUX2X1
XMUX2X1_38 MUX2X1_38/A MUX2X1_38/B XOR2X1_4/A gnd MUX2X1_57/A vdd MUX2X1
XMUX2X1_49 MUX2X1_49/A MUX2X1_49/B MUX2X1_49/S gnd MUX2X1_49/Y vdd MUX2X1
XINVX1_231 INVX1_231/A gnd INVX1_231/Y vdd INVX1
XINVX1_242 operand_B[59] gnd INVX1_242/Y vdd INVX1
XINVX1_253 INVX1_253/A gnd INVX1_253/Y vdd INVX1
XINVX1_275 BUFX2_29/A gnd INVX1_275/Y vdd INVX1
XINVX1_220 INVX1_220/A gnd INVX1_220/Y vdd INVX1
XINVX1_286 INVX1_286/A gnd INVX1_286/Y vdd INVX1
XINVX1_297 INVX1_297/A gnd INVX1_297/Y vdd INVX1
XINVX1_264 BUFX2_12/A gnd INVX1_264/Y vdd INVX1
XNAND2X1_97 BUFX4_69/Y OAI21X1_47/Y gnd OAI21X1_48/C vdd NAND2X1
XNAND2X1_53 operand_A[25] INVX1_23/Y gnd NAND2X1_55/A vdd NAND2X1
XNAND2X1_20 BUFX4_43/Y operand_A[0] gnd INVX2_10/A vdd NAND2X1
XNAND2X1_64 NOR2X1_48/Y OAI21X1_26/Y gnd NAND2X1_66/B vdd NAND2X1
XNAND2X1_75 XNOR2X1_4/Y XNOR2X1_5/Y gnd INVX1_82/A vdd NAND2X1
XNAND2X1_42 INVX2_27/Y INVX2_28/Y gnd NAND2X1_42/Y vdd NAND2X1
XNAND2X1_31 operand_A[14] INVX1_16/Y gnd INVX2_18/A vdd NAND2X1
XNAND2X1_86 MUX2X1_5/S operand_A[17] gnd OAI21X1_37/C vdd NAND2X1
XAOI21X1_246 NAND3X1_35/Y AOI21X1_246/B NOR2X1_336/Y gnd DFFPOSX1_60/D vdd AOI21X1
XAOI21X1_202 INVX1_224/Y INVX1_225/Y BUFX4_93/Y gnd AOI21X1_207/B vdd AOI21X1
XAOI21X1_257 OAI21X1_600/Y NOR2X1_352/Y NOR2X1_353/Y gnd DFFPOSX1_61/D vdd AOI21X1
XAOI21X1_224 INVX2_82/Y NOR2X1_321/Y BUFX4_30/Y gnd OAI21X1_572/C vdd AOI21X1
XAOI21X1_213 BUFX4_80/Y OAI22X1_33/B NAND3X1_33/Y gnd NAND2X1_485/A vdd AOI21X1
XAOI21X1_235 XOR2X1_7/A MUX2X1_51/B BUFX4_41/Y gnd AOI22X1_26/B vdd AOI21X1
XAOI21X1_268 INVX2_49/A INVX1_56/A INVX4_18/A gnd OAI21X1_625/C vdd AOI21X1
XAOI22X1_51 BUFX4_150/Y INVX1_321/Y BUFX4_3/Y AOI22X1_51/D gnd AOI22X1_51/Y vdd AOI22X1
XAOI21X1_279 XNOR2X1_18/Y INVX1_281/Y NOR2X1_21/Y gnd OAI21X1_644/C vdd AOI21X1
XAOI22X1_40 BUFX4_11/Y INVX1_263/Y AOI22X1_40/C AOI22X1_40/D gnd AOI22X1_40/Y vdd
+ AOI22X1
XOAI22X1_2 AND2X2_3/Y OAI22X1_2/B OAI22X1_2/C OAI22X1_2/D gnd OAI22X1_2/Y vdd OAI22X1
XNAND2X1_408 INVX4_14/Y INVX1_179/Y gnd NAND2X1_409/B vdd NAND2X1
XNAND2X1_419 BUFX4_38/Y NOR2X1_165/B gnd OAI21X1_446/C vdd NAND2X1
XNOR2X1_463 OR2X2_1/B AOI21X1_9/Y gnd NOR2X1_463/Y vdd NOR2X1
XNOR2X1_441 NOR2X1_441/A NOR2X1_441/B gnd NOR2X1_441/Y vdd NOR2X1
XNOR2X1_474 MUX2X1_57/S OAI22X1_1/A gnd NOR2X1_474/Y vdd NOR2X1
XNOR2X1_430 BUFX4_97/Y BUFX2_5/A gnd NOR2X1_430/Y vdd NOR2X1
XNOR2X1_452 BUFX4_82/Y NOR2X1_452/B gnd NOR2X1_452/Y vdd NOR2X1
XNOR2X1_485 NOR2X1_66/B NOR2X1_485/B gnd NOR2X1_486/B vdd NOR2X1
XOAI21X1_947 operand_B[29] operand_A[29] BUFX4_6/Y gnd OAI21X1_948/C vdd OAI21X1
XOAI21X1_936 BUFX4_158/Y XNOR2X1_26/Y BUFX4_99/Y gnd NOR2X1_503/A vdd OAI21X1
XOAI21X1_914 OAI21X1_23/A XNOR2X1_29/Y INVX1_323/Y gnd OAI21X1_915/A vdd OAI21X1
XOAI21X1_903 OAI21X1_903/A BUFX4_169/Y BUFX4_113/Y gnd OAI22X1_32/B vdd OAI21X1
XNOR2X1_496 NOR2X1_496/A OR2X2_49/A gnd NOR2X1_496/Y vdd NOR2X1
XOAI21X1_925 INVX1_324/Y BUFX4_167/Y OAI21X1_925/C gnd OAI21X1_925/Y vdd OAI21X1
XINVX2_44 operand_A[36] gnd INVX2_44/Y vdd INVX2
XINVX2_33 INVX2_33/A gnd INVX2_33/Y vdd INVX2
XINVX2_11 operand_A[3] gnd INVX2_11/Y vdd INVX2
XINVX2_22 operand_A[10] gnd INVX2_22/Y vdd INVX2
XINVX2_66 operand_A[38] gnd INVX2_66/Y vdd INVX2
XINVX2_77 operand_B[51] gnd INVX2_77/Y vdd INVX2
XINVX2_55 operand_A[37] gnd INVX2_55/Y vdd INVX2
XINVX2_88 INVX2_88/A gnd INVX2_88/Y vdd INVX2
XOAI21X1_29 OR2X2_3/A OAI21X1_29/B OAI21X1_29/C gnd OAI21X1_29/Y vdd OAI21X1
XOAI21X1_18 NOR2X1_29/B INVX1_312/A OAI21X1_18/C gnd OAI21X1_18/Y vdd OAI21X1
XNAND2X1_216 INVX8_1/A MUX2X1_8/Y gnd OAI21X1_183/C vdd NAND2X1
XNAND2X1_205 INVX1_31/Y NOR2X1_120/Y gnd OAI21X1_168/B vdd NAND2X1
XNAND2X1_249 NOR2X1_82/A OAI21X1_106/Y gnd OAI21X1_218/C vdd NAND2X1
XNAND2X1_238 INVX8_1/A MUX2X1_12/Y gnd OAI21X1_207/C vdd NAND2X1
XNAND2X1_227 BUFX4_67/Y INVX1_38/A gnd OAI21X1_194/C vdd NAND2X1
XNOR2X1_260 BUFX4_102/Y BUFX2_53/A gnd NOR2X1_260/Y vdd NOR2X1
XNOR2X1_293 operand_B[52] INVX2_40/Y gnd NOR2X1_293/Y vdd NOR2X1
XNOR2X1_271 INVX1_214/A NOR2X1_271/B gnd INVX1_212/A vdd NOR2X1
XNOR2X1_282 OAI22X1_11/Y OAI22X1_12/Y gnd NOR2X1_282/Y vdd NOR2X1
XOAI21X1_733 INVX1_294/Y XOR2X1_3/A OAI21X1_733/C gnd OAI21X1_734/B vdd OAI21X1
XOAI21X1_722 BUFX4_71/Y MUX2X1_70/Y OAI21X1_722/C gnd MUX2X1_111/A vdd OAI21X1
XOAI21X1_788 BUFX4_154/Y XNOR2X1_18/Y OAI21X1_788/C gnd NOR2X1_451/A vdd OAI21X1
XOAI21X1_744 XNOR2X1_17/Y OAI21X1_744/B OAI21X1_744/C gnd NAND3X1_59/B vdd OAI21X1
XOAI21X1_777 NOR2X1_448/Y OAI21X1_777/B OAI21X1_777/C gnd OAI21X1_777/Y vdd OAI21X1
XOAI21X1_700 XOR2X1_3/Y INVX2_10/Y NOR2X1_428/Y gnd OAI21X1_700/Y vdd OAI21X1
XOAI21X1_799 BUFX4_154/Y INVX1_17/A OAI21X1_799/C gnd NOR2X1_453/A vdd OAI21X1
XOAI21X1_755 BUFX4_62/Y OAI21X1_12/C BUFX4_97/Y gnd NOR2X1_440/A vdd OAI21X1
XOAI21X1_766 NAND3X1_62/Y NAND3X1_61/Y BUFX4_97/Y gnd OAI21X1_767/C vdd OAI21X1
XOAI21X1_711 INVX1_290/Y BUFX4_134/Y OAI21X1_711/C gnd MUX2X1_119/A vdd OAI21X1
XBUFX4_95 INVX8_11/Y gnd BUFX4_95/Y vdd BUFX4
XBUFX4_73 INVX8_1/Y gnd BUFX4_73/Y vdd BUFX4
XBUFX4_62 INVX8_17/Y gnd BUFX4_62/Y vdd BUFX4
XBUFX4_51 operand_B[0] gnd MUX2X1_6/S vdd BUFX4
XBUFX4_40 operand_B[3] gnd OR2X2_13/B vdd BUFX4
XBUFX4_84 BUFX4_87/A gnd BUFX4_84/Y vdd BUFX4
XOR2X2_21 OR2X2_21/A OR2X2_21/B gnd OR2X2_21/Y vdd OR2X2
XOR2X2_32 OR2X2_32/A OR2X2_32/B gnd OR2X2_32/Y vdd OR2X2
XOR2X2_10 OR2X2_10/A INVX8_5/A gnd OR2X2_10/Y vdd OR2X2
XXNOR2X1_5 operand_A[12] operand_B[12] gnd XNOR2X1_5/Y vdd XNOR2X1
XOR2X2_3 OR2X2_3/A OR2X2_3/B gnd OR2X2_3/Y vdd OR2X2
XOR2X2_43 OR2X2_43/A OR2X2_43/B gnd OR2X2_43/Y vdd OR2X2
XFILL_26_5_0 gnd vdd FILL
XFILL_1_5_0 gnd vdd FILL
XOAI21X1_530 BUFX4_102/Y INVX1_215/Y OAI21X1_530/C gnd OAI21X1_530/Y vdd OAI21X1
XINVX8_10 INVX8_10/A gnd INVX8_10/Y vdd INVX8
XOAI21X1_541 INVX1_138/A BUFX4_183/Y OAI21X1_541/C gnd OR2X2_32/A vdd OAI21X1
XINVX1_5 operand_B[17] gnd INVX1_5/Y vdd INVX1
XOAI21X1_552 OR2X2_33/B OAI21X1_552/B OAI21X1_552/C gnd OAI21X1_552/Y vdd OAI21X1
XOAI21X1_563 OAI21X1_563/A NOR2X1_307/A AND2X2_36/Y gnd OAI21X1_599/B vdd OAI21X1
XOAI21X1_596 INVX1_241/Y INVX1_244/A INVX1_243/Y gnd OAI21X1_596/Y vdd OAI21X1
XOAI21X1_585 OAI21X1_610/A INVX1_237/Y INVX1_240/Y gnd AND2X2_41/A vdd OAI21X1
XOAI21X1_574 NOR2X1_320/B NOR2X1_320/A NOR2X1_323/A gnd OAI21X1_584/C vdd OAI21X1
.ends

